`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/05/24 09:32:12
// Design Name: 
// Module Name: cnn
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cnn(
clk, rst_n, Start, ReadEn
    );
    input clk;
    input rst_n;
    input Start;
    input ReadEn;
    
    
    reg   [7:0]   Image   [1023:0];
    reg   [35:0]  Filter = 36'b000100010001000110010001000100010001;
    reg   [15:0]    Conv_out    [899:0];
//    reg   [7:0]   Filter  [8:0];
    reg   [35:0]    Filter_0 = 36'b000100010001000110010001000100010001;
    reg   [31:0]    Conv_out_2    [783:0];
    initial begin 
    $readmemh("input.mem", Image);
//    $readmemh("filter.mem", Filter);
    end
    wire    [71:0]  image_0_0, image_0_1, image_0_2, image_0_3, image_0_4, image_0_5, image_0_6, image_0_7, image_0_8, image_0_9;
    wire    [71:0]  image_0_10, image_0_11, image_0_12, image_0_13, image_0_14, image_0_15, image_0_16, image_0_17, image_0_18, image_0_19;
    wire    [71:0]  image_0_20, image_0_21, image_0_22, image_0_23, image_0_24, image_0_25, image_0_26, image_0_27, image_0_28, image_0_29;
    wire    [71:0]  image_0_30, image_0_31, image_0_32, image_0_33, image_0_34, image_0_35, image_0_36, image_0_37, image_0_38, image_0_39;
    wire    [71:0]  image_0_40, image_0_41, image_0_42, image_0_43, image_0_44, image_0_45, image_0_46, image_0_47, image_0_48, image_0_49;
    wire    [71:0]  image_0_50, image_0_51, image_0_52, image_0_53, image_0_54, image_0_55, image_0_56, image_0_57, image_0_58, image_0_59;
    wire    [71:0]  image_0_60, image_0_61, image_0_62, image_0_63, image_0_64, image_0_65, image_0_66, image_0_67, image_0_68, image_0_69;
    wire    [71:0]  image_0_70, image_0_71, image_0_72, image_0_73, image_0_74, image_0_75, image_0_76, image_0_77, image_0_78, image_0_79;
    wire    [71:0]  image_0_80, image_0_81, image_0_82, image_0_83, image_0_84, image_0_85, image_0_86, image_0_87, image_0_88, image_0_89;
    wire    [71:0]  image_0_90, image_0_91, image_0_92, image_0_93, image_0_94, image_0_95, image_0_96, image_0_97, image_0_98, image_0_99;
    wire    [71:0]  image_0_100, image_0_101, image_0_102, image_0_103, image_0_104, image_0_105, image_0_106, image_0_107, image_0_108, image_0_109;
    wire    [71:0]  image_0_110, image_0_111, image_0_112, image_0_113, image_0_114, image_0_115, image_0_116, image_0_117, image_0_118, image_0_119;
    wire    [71:0]  image_0_120, image_0_121, image_0_122, image_0_123, image_0_124, image_0_125, image_0_126, image_0_127, image_0_128, image_0_129;
    wire    [71:0]  image_0_130, image_0_131, image_0_132, image_0_133, image_0_134, image_0_135, image_0_136, image_0_137, image_0_138, image_0_139;
    wire    [71:0]  image_0_140, image_0_141, image_0_142, image_0_143, image_0_144, image_0_145, image_0_146, image_0_147, image_0_148, image_0_149;
    wire    [71:0]  image_0_150, image_0_151, image_0_152, image_0_153, image_0_154, image_0_155, image_0_156, image_0_157, image_0_158, image_0_159;
    wire    [71:0]  image_0_160, image_0_161, image_0_162, image_0_163, image_0_164, image_0_165, image_0_166, image_0_167, image_0_168, image_0_169;
    wire    [71:0]  image_0_170, image_0_171, image_0_172, image_0_173, image_0_174, image_0_175, image_0_176, image_0_177, image_0_178, image_0_179;
    wire    [71:0]  image_0_180, image_0_181, image_0_182, image_0_183, image_0_184, image_0_185, image_0_186, image_0_187, image_0_188, image_0_189;
    wire    [71:0]  image_0_190, image_0_191, image_0_192, image_0_193, image_0_194, image_0_195, image_0_196, image_0_197, image_0_198, image_0_199;
    wire    [71:0]  image_0_200, image_0_201, image_0_202, image_0_203, image_0_204, image_0_205, image_0_206, image_0_207, image_0_208, image_0_209;
    wire    [71:0]  image_0_210, image_0_211, image_0_212, image_0_213, image_0_214, image_0_215, image_0_216, image_0_217, image_0_218, image_0_219;
    wire    [71:0]  image_0_220, image_0_221, image_0_222, image_0_223, image_0_224, image_0_225, image_0_226, image_0_227, image_0_228, image_0_229;
    wire    [71:0]  image_0_230, image_0_231, image_0_232, image_0_233, image_0_234, image_0_235, image_0_236, image_0_237, image_0_238, image_0_239;
    wire    [71:0]  image_0_240, image_0_241, image_0_242, image_0_243, image_0_244, image_0_245, image_0_246, image_0_247, image_0_248, image_0_249;
    wire    [71:0]  image_0_250, image_0_251, image_0_252, image_0_253, image_0_254, image_0_255, image_0_256, image_0_257, image_0_258, image_0_259;
    wire    [71:0]  image_0_260, image_0_261, image_0_262, image_0_263, image_0_264, image_0_265, image_0_266, image_0_267, image_0_268, image_0_269;
    wire    [71:0]  image_0_270, image_0_271, image_0_272, image_0_273, image_0_274, image_0_275, image_0_276, image_0_277, image_0_278, image_0_279;
    wire    [71:0]  image_0_280, image_0_281, image_0_282, image_0_283, image_0_284, image_0_285, image_0_286, image_0_287, image_0_288, image_0_289;
    wire    [71:0]  image_0_290, image_0_291, image_0_292, image_0_293, image_0_294, image_0_295, image_0_296, image_0_297, image_0_298, image_0_299;
    wire    [71:0]  image_0_300, image_0_301, image_0_302, image_0_303, image_0_304, image_0_305, image_0_306, image_0_307, image_0_308, image_0_309;
    wire    [71:0]  image_0_310, image_0_311, image_0_312, image_0_313, image_0_314, image_0_315, image_0_316, image_0_317, image_0_318, image_0_319;
    wire    [71:0]  image_0_320, image_0_321, image_0_322, image_0_323, image_0_324, image_0_325, image_0_326, image_0_327, image_0_328, image_0_329;
    wire    [71:0]  image_0_330, image_0_331, image_0_332, image_0_333, image_0_334, image_0_335, image_0_336, image_0_337, image_0_338, image_0_339;
    wire    [71:0]  image_0_340, image_0_341, image_0_342, image_0_343, image_0_344, image_0_345, image_0_346, image_0_347, image_0_348, image_0_349;
    wire    [71:0]  image_0_350, image_0_351, image_0_352, image_0_353, image_0_354, image_0_355, image_0_356, image_0_357, image_0_358, image_0_359;
    wire    [71:0]  image_0_360, image_0_361, image_0_362, image_0_363, image_0_364, image_0_365, image_0_366, image_0_367, image_0_368, image_0_369;
    wire    [71:0]  image_0_370, image_0_371, image_0_372, image_0_373, image_0_374, image_0_375, image_0_376, image_0_377, image_0_378, image_0_379;
    wire    [71:0]  image_0_380, image_0_381, image_0_382, image_0_383, image_0_384, image_0_385, image_0_386, image_0_387, image_0_388, image_0_389;
    wire    [71:0]  image_0_390, image_0_391, image_0_392, image_0_393, image_0_394, image_0_395, image_0_396, image_0_397, image_0_398, image_0_399;
    wire    [71:0]  image_0_400, image_0_401, image_0_402, image_0_403, image_0_404, image_0_405, image_0_406, image_0_407, image_0_408, image_0_409;
    wire    [71:0]  image_0_410, image_0_411, image_0_412, image_0_413, image_0_414, image_0_415, image_0_416, image_0_417, image_0_418, image_0_419;
    wire    [71:0]  image_0_420, image_0_421, image_0_422, image_0_423, image_0_424, image_0_425, image_0_426, image_0_427, image_0_428, image_0_429;
    wire    [71:0]  image_0_430, image_0_431, image_0_432, image_0_433, image_0_434, image_0_435, image_0_436, image_0_437, image_0_438, image_0_439;
    wire    [71:0]  image_0_440, image_0_441, image_0_442, image_0_443, image_0_444, image_0_445, image_0_446, image_0_447, image_0_448, image_0_449;
    wire    [71:0]  image_0_450, image_0_451, image_0_452, image_0_453, image_0_454, image_0_455, image_0_456, image_0_457, image_0_458, image_0_459;
    wire    [71:0]  image_0_460, image_0_461, image_0_462, image_0_463, image_0_464, image_0_465, image_0_466, image_0_467, image_0_468, image_0_469;
    wire    [71:0]  image_0_470, image_0_471, image_0_472, image_0_473, image_0_474, image_0_475, image_0_476, image_0_477, image_0_478, image_0_479;
    wire    [71:0]  image_0_480, image_0_481, image_0_482, image_0_483, image_0_484, image_0_485, image_0_486, image_0_487, image_0_488, image_0_489;
    wire    [71:0]  image_0_490, image_0_491, image_0_492, image_0_493, image_0_494, image_0_495, image_0_496, image_0_497, image_0_498, image_0_499;
    wire    [71:0]  image_0_500, image_0_501, image_0_502, image_0_503, image_0_504, image_0_505, image_0_506, image_0_507, image_0_508, image_0_509;
    wire    [71:0]  image_0_510, image_0_511, image_0_512, image_0_513, image_0_514, image_0_515, image_0_516, image_0_517, image_0_518, image_0_519;
    wire    [71:0]  image_0_520, image_0_521, image_0_522, image_0_523, image_0_524, image_0_525, image_0_526, image_0_527, image_0_528, image_0_529;
    wire    [71:0]  image_0_530, image_0_531, image_0_532, image_0_533, image_0_534, image_0_535, image_0_536, image_0_537, image_0_538, image_0_539;
    wire    [71:0]  image_0_540, image_0_541, image_0_542, image_0_543, image_0_544, image_0_545, image_0_546, image_0_547, image_0_548, image_0_549;
    wire    [71:0]  image_0_550, image_0_551, image_0_552, image_0_553, image_0_554, image_0_555, image_0_556, image_0_557, image_0_558, image_0_559;
    wire    [71:0]  image_0_560, image_0_561, image_0_562, image_0_563, image_0_564, image_0_565, image_0_566, image_0_567, image_0_568, image_0_569;
    wire    [71:0]  image_0_570, image_0_571, image_0_572, image_0_573, image_0_574, image_0_575, image_0_576, image_0_577, image_0_578, image_0_579;
    wire    [71:0]  image_0_580, image_0_581, image_0_582, image_0_583, image_0_584, image_0_585, image_0_586, image_0_587, image_0_588, image_0_589;
    wire    [71:0]  image_0_590, image_0_591, image_0_592, image_0_593, image_0_594, image_0_595, image_0_596, image_0_597, image_0_598, image_0_599;
    wire    [71:0]  image_0_600, image_0_601, image_0_602, image_0_603, image_0_604, image_0_605, image_0_606, image_0_607, image_0_608, image_0_609;
    wire    [71:0]  image_0_610, image_0_611, image_0_612, image_0_613, image_0_614, image_0_615, image_0_616, image_0_617, image_0_618, image_0_619;
    wire    [71:0]  image_0_620, image_0_621, image_0_622, image_0_623, image_0_624, image_0_625, image_0_626, image_0_627, image_0_628, image_0_629;
    wire    [71:0]  image_0_630, image_0_631, image_0_632, image_0_633, image_0_634, image_0_635, image_0_636, image_0_637, image_0_638, image_0_639;
    wire    [71:0]  image_0_640, image_0_641, image_0_642, image_0_643, image_0_644, image_0_645, image_0_646, image_0_647, image_0_648, image_0_649;
    wire    [71:0]  image_0_650, image_0_651, image_0_652, image_0_653, image_0_654, image_0_655, image_0_656, image_0_657, image_0_658, image_0_659;
    wire    [71:0]  image_0_660, image_0_661, image_0_662, image_0_663, image_0_664, image_0_665, image_0_666, image_0_667, image_0_668, image_0_669;
    wire    [71:0]  image_0_670, image_0_671, image_0_672, image_0_673, image_0_674, image_0_675, image_0_676, image_0_677, image_0_678, image_0_679;
    wire    [71:0]  image_0_680, image_0_681, image_0_682, image_0_683, image_0_684, image_0_685, image_0_686, image_0_687, image_0_688, image_0_689;
    wire    [71:0]  image_0_690, image_0_691, image_0_692, image_0_693, image_0_694, image_0_695, image_0_696, image_0_697, image_0_698, image_0_699;
    wire    [71:0]  image_0_700, image_0_701, image_0_702, image_0_703, image_0_704, image_0_705, image_0_706, image_0_707, image_0_708, image_0_709;
    wire    [71:0]  image_0_710, image_0_711, image_0_712, image_0_713, image_0_714, image_0_715, image_0_716, image_0_717, image_0_718, image_0_719;
    wire    [71:0]  image_0_720, image_0_721, image_0_722, image_0_723, image_0_724, image_0_725, image_0_726, image_0_727, image_0_728, image_0_729;
    wire    [71:0]  image_0_730, image_0_731, image_0_732, image_0_733, image_0_734, image_0_735, image_0_736, image_0_737, image_0_738, image_0_739;
    wire    [71:0]  image_0_740, image_0_741, image_0_742, image_0_743, image_0_744, image_0_745, image_0_746, image_0_747, image_0_748, image_0_749;
    wire    [71:0]  image_0_750, image_0_751, image_0_752, image_0_753, image_0_754, image_0_755, image_0_756, image_0_757, image_0_758, image_0_759;
    wire    [71:0]  image_0_760, image_0_761, image_0_762, image_0_763, image_0_764, image_0_765, image_0_766, image_0_767, image_0_768, image_0_769;
    wire    [71:0]  image_0_770, image_0_771, image_0_772, image_0_773, image_0_774, image_0_775, image_0_776, image_0_777, image_0_778, image_0_779;
    wire    [71:0]  image_0_780, image_0_781, image_0_782, image_0_783, image_0_784, image_0_785, image_0_786, image_0_787, image_0_788, image_0_789;
    wire    [71:0]  image_0_790, image_0_791, image_0_792, image_0_793, image_0_794, image_0_795, image_0_796, image_0_797, image_0_798, image_0_799;
    wire    [71:0]  image_0_800, image_0_801, image_0_802, image_0_803, image_0_804, image_0_805, image_0_806, image_0_807, image_0_808, image_0_809;
    wire    [71:0]  image_0_810, image_0_811, image_0_812, image_0_813, image_0_814, image_0_815, image_0_816, image_0_817, image_0_818, image_0_819;
    wire    [71:0]  image_0_820, image_0_821, image_0_822, image_0_823, image_0_824, image_0_825, image_0_826, image_0_827, image_0_828, image_0_829;
    wire    [71:0]  image_0_830, image_0_831, image_0_832, image_0_833, image_0_834, image_0_835, image_0_836, image_0_837, image_0_838, image_0_839;
    wire    [71:0]  image_0_840, image_0_841, image_0_842, image_0_843, image_0_844, image_0_845, image_0_846, image_0_847, image_0_848, image_0_849;
    wire    [71:0]  image_0_850, image_0_851, image_0_852, image_0_853, image_0_854, image_0_855, image_0_856, image_0_857, image_0_858, image_0_859;
    wire    [71:0]  image_0_860, image_0_861, image_0_862, image_0_863, image_0_864, image_0_865, image_0_866, image_0_867, image_0_868, image_0_869;
    wire    [71:0]  image_0_870, image_0_871, image_0_872, image_0_873, image_0_874, image_0_875, image_0_876, image_0_877, image_0_878, image_0_879;
    wire    [71:0]  image_0_880, image_0_881, image_0_882, image_0_883, image_0_884, image_0_885, image_0_886, image_0_887, image_0_888, image_0_889;
    wire    [71:0]  image_0_890, image_0_891, image_0_892, image_0_893, image_0_894, image_0_895, image_0_896, image_0_897, image_0_898, image_0_899;

wire    [15:0]  conv_out_0_0, conv_out_0_1, conv_out_0_2, conv_out_0_3, conv_out_0_4, conv_out_0_5, conv_out_0_6, conv_out_0_7, conv_out_0_8, conv_out_0_9;
wire    [15:0]  conv_out_0_10, conv_out_0_11, conv_out_0_12, conv_out_0_13, conv_out_0_14, conv_out_0_15, conv_out_0_16, conv_out_0_17, conv_out_0_18, conv_out_0_19;
wire    [15:0]  conv_out_0_20, conv_out_0_21, conv_out_0_22, conv_out_0_23, conv_out_0_24, conv_out_0_25, conv_out_0_26, conv_out_0_27, conv_out_0_28, conv_out_0_29;
wire    [15:0]  conv_out_0_30, conv_out_0_31, conv_out_0_32, conv_out_0_33, conv_out_0_34, conv_out_0_35, conv_out_0_36, conv_out_0_37, conv_out_0_38, conv_out_0_39;
wire    [15:0]  conv_out_0_40, conv_out_0_41, conv_out_0_42, conv_out_0_43, conv_out_0_44, conv_out_0_45, conv_out_0_46, conv_out_0_47, conv_out_0_48, conv_out_0_49;
wire    [15:0]  conv_out_0_50, conv_out_0_51, conv_out_0_52, conv_out_0_53, conv_out_0_54, conv_out_0_55, conv_out_0_56, conv_out_0_57, conv_out_0_58, conv_out_0_59;
wire    [15:0]  conv_out_0_60, conv_out_0_61, conv_out_0_62, conv_out_0_63, conv_out_0_64, conv_out_0_65, conv_out_0_66, conv_out_0_67, conv_out_0_68, conv_out_0_69;
wire    [15:0]  conv_out_0_70, conv_out_0_71, conv_out_0_72, conv_out_0_73, conv_out_0_74, conv_out_0_75, conv_out_0_76, conv_out_0_77, conv_out_0_78, conv_out_0_79;
wire    [15:0]  conv_out_0_80, conv_out_0_81, conv_out_0_82, conv_out_0_83, conv_out_0_84, conv_out_0_85, conv_out_0_86, conv_out_0_87, conv_out_0_88, conv_out_0_89;
wire    [15:0]  conv_out_0_90, conv_out_0_91, conv_out_0_92, conv_out_0_93, conv_out_0_94, conv_out_0_95, conv_out_0_96, conv_out_0_97, conv_out_0_98, conv_out_0_99;
wire    [15:0]  conv_out_0_100, conv_out_0_101, conv_out_0_102, conv_out_0_103, conv_out_0_104, conv_out_0_105, conv_out_0_106, conv_out_0_107, conv_out_0_108, conv_out_0_109;
wire    [15:0]  conv_out_0_110, conv_out_0_111, conv_out_0_112, conv_out_0_113, conv_out_0_114, conv_out_0_115, conv_out_0_116, conv_out_0_117, conv_out_0_118, conv_out_0_119;
wire    [15:0]  conv_out_0_120, conv_out_0_121, conv_out_0_122, conv_out_0_123, conv_out_0_124, conv_out_0_125, conv_out_0_126, conv_out_0_127, conv_out_0_128, conv_out_0_129;
wire    [15:0]  conv_out_0_130, conv_out_0_131, conv_out_0_132, conv_out_0_133, conv_out_0_134, conv_out_0_135, conv_out_0_136, conv_out_0_137, conv_out_0_138, conv_out_0_139;
wire    [15:0]  conv_out_0_140, conv_out_0_141, conv_out_0_142, conv_out_0_143, conv_out_0_144, conv_out_0_145, conv_out_0_146, conv_out_0_147, conv_out_0_148, conv_out_0_149;
wire    [15:0]  conv_out_0_150, conv_out_0_151, conv_out_0_152, conv_out_0_153, conv_out_0_154, conv_out_0_155, conv_out_0_156, conv_out_0_157, conv_out_0_158, conv_out_0_159;
wire    [15:0]  conv_out_0_160, conv_out_0_161, conv_out_0_162, conv_out_0_163, conv_out_0_164, conv_out_0_165, conv_out_0_166, conv_out_0_167, conv_out_0_168, conv_out_0_169;
wire    [15:0]  conv_out_0_170, conv_out_0_171, conv_out_0_172, conv_out_0_173, conv_out_0_174, conv_out_0_175, conv_out_0_176, conv_out_0_177, conv_out_0_178, conv_out_0_179;
wire    [15:0]  conv_out_0_180, conv_out_0_181, conv_out_0_182, conv_out_0_183, conv_out_0_184, conv_out_0_185, conv_out_0_186, conv_out_0_187, conv_out_0_188, conv_out_0_189;
wire    [15:0]  conv_out_0_190, conv_out_0_191, conv_out_0_192, conv_out_0_193, conv_out_0_194, conv_out_0_195, conv_out_0_196, conv_out_0_197, conv_out_0_198, conv_out_0_199;
wire    [15:0]  conv_out_0_200, conv_out_0_201, conv_out_0_202, conv_out_0_203, conv_out_0_204, conv_out_0_205, conv_out_0_206, conv_out_0_207, conv_out_0_208, conv_out_0_209;
wire    [15:0]  conv_out_0_210, conv_out_0_211, conv_out_0_212, conv_out_0_213, conv_out_0_214, conv_out_0_215, conv_out_0_216, conv_out_0_217, conv_out_0_218, conv_out_0_219;
wire    [15:0]  conv_out_0_220, conv_out_0_221, conv_out_0_222, conv_out_0_223, conv_out_0_224, conv_out_0_225, conv_out_0_226, conv_out_0_227, conv_out_0_228, conv_out_0_229;
wire    [15:0]  conv_out_0_230, conv_out_0_231, conv_out_0_232, conv_out_0_233, conv_out_0_234, conv_out_0_235, conv_out_0_236, conv_out_0_237, conv_out_0_238, conv_out_0_239;
wire    [15:0]  conv_out_0_240, conv_out_0_241, conv_out_0_242, conv_out_0_243, conv_out_0_244, conv_out_0_245, conv_out_0_246, conv_out_0_247, conv_out_0_248, conv_out_0_249;
wire    [15:0]  conv_out_0_250, conv_out_0_251, conv_out_0_252, conv_out_0_253, conv_out_0_254, conv_out_0_255, conv_out_0_256, conv_out_0_257, conv_out_0_258, conv_out_0_259;
wire    [15:0]  conv_out_0_260, conv_out_0_261, conv_out_0_262, conv_out_0_263, conv_out_0_264, conv_out_0_265, conv_out_0_266, conv_out_0_267, conv_out_0_268, conv_out_0_269;
wire    [15:0]  conv_out_0_270, conv_out_0_271, conv_out_0_272, conv_out_0_273, conv_out_0_274, conv_out_0_275, conv_out_0_276, conv_out_0_277, conv_out_0_278, conv_out_0_279;
wire    [15:0]  conv_out_0_280, conv_out_0_281, conv_out_0_282, conv_out_0_283, conv_out_0_284, conv_out_0_285, conv_out_0_286, conv_out_0_287, conv_out_0_288, conv_out_0_289;
wire    [15:0]  conv_out_0_290, conv_out_0_291, conv_out_0_292, conv_out_0_293, conv_out_0_294, conv_out_0_295, conv_out_0_296, conv_out_0_297, conv_out_0_298, conv_out_0_299;
wire    [15:0]  conv_out_0_300, conv_out_0_301, conv_out_0_302, conv_out_0_303, conv_out_0_304, conv_out_0_305, conv_out_0_306, conv_out_0_307, conv_out_0_308, conv_out_0_309;
wire    [15:0]  conv_out_0_310, conv_out_0_311, conv_out_0_312, conv_out_0_313, conv_out_0_314, conv_out_0_315, conv_out_0_316, conv_out_0_317, conv_out_0_318, conv_out_0_319;
wire    [15:0]  conv_out_0_320, conv_out_0_321, conv_out_0_322, conv_out_0_323, conv_out_0_324, conv_out_0_325, conv_out_0_326, conv_out_0_327, conv_out_0_328, conv_out_0_329;
wire    [15:0]  conv_out_0_330, conv_out_0_331, conv_out_0_332, conv_out_0_333, conv_out_0_334, conv_out_0_335, conv_out_0_336, conv_out_0_337, conv_out_0_338, conv_out_0_339;
wire    [15:0]  conv_out_0_340, conv_out_0_341, conv_out_0_342, conv_out_0_343, conv_out_0_344, conv_out_0_345, conv_out_0_346, conv_out_0_347, conv_out_0_348, conv_out_0_349;
wire    [15:0]  conv_out_0_350, conv_out_0_351, conv_out_0_352, conv_out_0_353, conv_out_0_354, conv_out_0_355, conv_out_0_356, conv_out_0_357, conv_out_0_358, conv_out_0_359;
wire    [15:0]  conv_out_0_360, conv_out_0_361, conv_out_0_362, conv_out_0_363, conv_out_0_364, conv_out_0_365, conv_out_0_366, conv_out_0_367, conv_out_0_368, conv_out_0_369;
wire    [15:0]  conv_out_0_370, conv_out_0_371, conv_out_0_372, conv_out_0_373, conv_out_0_374, conv_out_0_375, conv_out_0_376, conv_out_0_377, conv_out_0_378, conv_out_0_379;
wire    [15:0]  conv_out_0_380, conv_out_0_381, conv_out_0_382, conv_out_0_383, conv_out_0_384, conv_out_0_385, conv_out_0_386, conv_out_0_387, conv_out_0_388, conv_out_0_389;
wire    [15:0]  conv_out_0_390, conv_out_0_391, conv_out_0_392, conv_out_0_393, conv_out_0_394, conv_out_0_395, conv_out_0_396, conv_out_0_397, conv_out_0_398, conv_out_0_399;
wire    [15:0]  conv_out_0_400, conv_out_0_401, conv_out_0_402, conv_out_0_403, conv_out_0_404, conv_out_0_405, conv_out_0_406, conv_out_0_407, conv_out_0_408, conv_out_0_409;
wire    [15:0]  conv_out_0_410, conv_out_0_411, conv_out_0_412, conv_out_0_413, conv_out_0_414, conv_out_0_415, conv_out_0_416, conv_out_0_417, conv_out_0_418, conv_out_0_419;
wire    [15:0]  conv_out_0_420, conv_out_0_421, conv_out_0_422, conv_out_0_423, conv_out_0_424, conv_out_0_425, conv_out_0_426, conv_out_0_427, conv_out_0_428, conv_out_0_429;
wire    [15:0]  conv_out_0_430, conv_out_0_431, conv_out_0_432, conv_out_0_433, conv_out_0_434, conv_out_0_435, conv_out_0_436, conv_out_0_437, conv_out_0_438, conv_out_0_439;
wire    [15:0]  conv_out_0_440, conv_out_0_441, conv_out_0_442, conv_out_0_443, conv_out_0_444, conv_out_0_445, conv_out_0_446, conv_out_0_447, conv_out_0_448, conv_out_0_449;
wire    [15:0]  conv_out_0_450, conv_out_0_451, conv_out_0_452, conv_out_0_453, conv_out_0_454, conv_out_0_455, conv_out_0_456, conv_out_0_457, conv_out_0_458, conv_out_0_459;
wire    [15:0]  conv_out_0_460, conv_out_0_461, conv_out_0_462, conv_out_0_463, conv_out_0_464, conv_out_0_465, conv_out_0_466, conv_out_0_467, conv_out_0_468, conv_out_0_469;
wire    [15:0]  conv_out_0_470, conv_out_0_471, conv_out_0_472, conv_out_0_473, conv_out_0_474, conv_out_0_475, conv_out_0_476, conv_out_0_477, conv_out_0_478, conv_out_0_479;
wire    [15:0]  conv_out_0_480, conv_out_0_481, conv_out_0_482, conv_out_0_483, conv_out_0_484, conv_out_0_485, conv_out_0_486, conv_out_0_487, conv_out_0_488, conv_out_0_489;
wire    [15:0]  conv_out_0_490, conv_out_0_491, conv_out_0_492, conv_out_0_493, conv_out_0_494, conv_out_0_495, conv_out_0_496, conv_out_0_497, conv_out_0_498, conv_out_0_499;
wire    [15:0]  conv_out_0_500, conv_out_0_501, conv_out_0_502, conv_out_0_503, conv_out_0_504, conv_out_0_505, conv_out_0_506, conv_out_0_507, conv_out_0_508, conv_out_0_509;
wire    [15:0]  conv_out_0_510, conv_out_0_511, conv_out_0_512, conv_out_0_513, conv_out_0_514, conv_out_0_515, conv_out_0_516, conv_out_0_517, conv_out_0_518, conv_out_0_519;
wire    [15:0]  conv_out_0_520, conv_out_0_521, conv_out_0_522, conv_out_0_523, conv_out_0_524, conv_out_0_525, conv_out_0_526, conv_out_0_527, conv_out_0_528, conv_out_0_529;
wire    [15:0]  conv_out_0_530, conv_out_0_531, conv_out_0_532, conv_out_0_533, conv_out_0_534, conv_out_0_535, conv_out_0_536, conv_out_0_537, conv_out_0_538, conv_out_0_539;
wire    [15:0]  conv_out_0_540, conv_out_0_541, conv_out_0_542, conv_out_0_543, conv_out_0_544, conv_out_0_545, conv_out_0_546, conv_out_0_547, conv_out_0_548, conv_out_0_549;
wire    [15:0]  conv_out_0_550, conv_out_0_551, conv_out_0_552, conv_out_0_553, conv_out_0_554, conv_out_0_555, conv_out_0_556, conv_out_0_557, conv_out_0_558, conv_out_0_559;
wire    [15:0]  conv_out_0_560, conv_out_0_561, conv_out_0_562, conv_out_0_563, conv_out_0_564, conv_out_0_565, conv_out_0_566, conv_out_0_567, conv_out_0_568, conv_out_0_569;
wire    [15:0]  conv_out_0_570, conv_out_0_571, conv_out_0_572, conv_out_0_573, conv_out_0_574, conv_out_0_575, conv_out_0_576, conv_out_0_577, conv_out_0_578, conv_out_0_579;
wire    [15:0]  conv_out_0_580, conv_out_0_581, conv_out_0_582, conv_out_0_583, conv_out_0_584, conv_out_0_585, conv_out_0_586, conv_out_0_587, conv_out_0_588, conv_out_0_589;
wire    [15:0]  conv_out_0_590, conv_out_0_591, conv_out_0_592, conv_out_0_593, conv_out_0_594, conv_out_0_595, conv_out_0_596, conv_out_0_597, conv_out_0_598, conv_out_0_599;
wire    [15:0]  conv_out_0_600, conv_out_0_601, conv_out_0_602, conv_out_0_603, conv_out_0_604, conv_out_0_605, conv_out_0_606, conv_out_0_607, conv_out_0_608, conv_out_0_609;
wire    [15:0]  conv_out_0_610, conv_out_0_611, conv_out_0_612, conv_out_0_613, conv_out_0_614, conv_out_0_615, conv_out_0_616, conv_out_0_617, conv_out_0_618, conv_out_0_619;
wire    [15:0]  conv_out_0_620, conv_out_0_621, conv_out_0_622, conv_out_0_623, conv_out_0_624, conv_out_0_625, conv_out_0_626, conv_out_0_627, conv_out_0_628, conv_out_0_629;
wire    [15:0]  conv_out_0_630, conv_out_0_631, conv_out_0_632, conv_out_0_633, conv_out_0_634, conv_out_0_635, conv_out_0_636, conv_out_0_637, conv_out_0_638, conv_out_0_639;
wire    [15:0]  conv_out_0_640, conv_out_0_641, conv_out_0_642, conv_out_0_643, conv_out_0_644, conv_out_0_645, conv_out_0_646, conv_out_0_647, conv_out_0_648, conv_out_0_649;
wire    [15:0]  conv_out_0_650, conv_out_0_651, conv_out_0_652, conv_out_0_653, conv_out_0_654, conv_out_0_655, conv_out_0_656, conv_out_0_657, conv_out_0_658, conv_out_0_659;
wire    [15:0]  conv_out_0_660, conv_out_0_661, conv_out_0_662, conv_out_0_663, conv_out_0_664, conv_out_0_665, conv_out_0_666, conv_out_0_667, conv_out_0_668, conv_out_0_669;
wire    [15:0]  conv_out_0_670, conv_out_0_671, conv_out_0_672, conv_out_0_673, conv_out_0_674, conv_out_0_675, conv_out_0_676, conv_out_0_677, conv_out_0_678, conv_out_0_679;
wire    [15:0]  conv_out_0_680, conv_out_0_681, conv_out_0_682, conv_out_0_683, conv_out_0_684, conv_out_0_685, conv_out_0_686, conv_out_0_687, conv_out_0_688, conv_out_0_689;
wire    [15:0]  conv_out_0_690, conv_out_0_691, conv_out_0_692, conv_out_0_693, conv_out_0_694, conv_out_0_695, conv_out_0_696, conv_out_0_697, conv_out_0_698, conv_out_0_699;
wire    [15:0]  conv_out_0_700, conv_out_0_701, conv_out_0_702, conv_out_0_703, conv_out_0_704, conv_out_0_705, conv_out_0_706, conv_out_0_707, conv_out_0_708, conv_out_0_709;
wire    [15:0]  conv_out_0_710, conv_out_0_711, conv_out_0_712, conv_out_0_713, conv_out_0_714, conv_out_0_715, conv_out_0_716, conv_out_0_717, conv_out_0_718, conv_out_0_719;
wire    [15:0]  conv_out_0_720, conv_out_0_721, conv_out_0_722, conv_out_0_723, conv_out_0_724, conv_out_0_725, conv_out_0_726, conv_out_0_727, conv_out_0_728, conv_out_0_729;
wire    [15:0]  conv_out_0_730, conv_out_0_731, conv_out_0_732, conv_out_0_733, conv_out_0_734, conv_out_0_735, conv_out_0_736, conv_out_0_737, conv_out_0_738, conv_out_0_739;
wire    [15:0]  conv_out_0_740, conv_out_0_741, conv_out_0_742, conv_out_0_743, conv_out_0_744, conv_out_0_745, conv_out_0_746, conv_out_0_747, conv_out_0_748, conv_out_0_749;
wire    [15:0]  conv_out_0_750, conv_out_0_751, conv_out_0_752, conv_out_0_753, conv_out_0_754, conv_out_0_755, conv_out_0_756, conv_out_0_757, conv_out_0_758, conv_out_0_759;
wire    [15:0]  conv_out_0_760, conv_out_0_761, conv_out_0_762, conv_out_0_763, conv_out_0_764, conv_out_0_765, conv_out_0_766, conv_out_0_767, conv_out_0_768, conv_out_0_769;
wire    [15:0]  conv_out_0_770, conv_out_0_771, conv_out_0_772, conv_out_0_773, conv_out_0_774, conv_out_0_775, conv_out_0_776, conv_out_0_777, conv_out_0_778, conv_out_0_779;
wire    [15:0]  conv_out_0_780, conv_out_0_781, conv_out_0_782, conv_out_0_783, conv_out_0_784, conv_out_0_785, conv_out_0_786, conv_out_0_787, conv_out_0_788, conv_out_0_789;
wire    [15:0]  conv_out_0_790, conv_out_0_791, conv_out_0_792, conv_out_0_793, conv_out_0_794, conv_out_0_795, conv_out_0_796, conv_out_0_797, conv_out_0_798, conv_out_0_799;
wire    [15:0]  conv_out_0_800, conv_out_0_801, conv_out_0_802, conv_out_0_803, conv_out_0_804, conv_out_0_805, conv_out_0_806, conv_out_0_807, conv_out_0_808, conv_out_0_809;
wire    [15:0]  conv_out_0_810, conv_out_0_811, conv_out_0_812, conv_out_0_813, conv_out_0_814, conv_out_0_815, conv_out_0_816, conv_out_0_817, conv_out_0_818, conv_out_0_819;
wire    [15:0]  conv_out_0_820, conv_out_0_821, conv_out_0_822, conv_out_0_823, conv_out_0_824, conv_out_0_825, conv_out_0_826, conv_out_0_827, conv_out_0_828, conv_out_0_829;
wire    [15:0]  conv_out_0_830, conv_out_0_831, conv_out_0_832, conv_out_0_833, conv_out_0_834, conv_out_0_835, conv_out_0_836, conv_out_0_837, conv_out_0_838, conv_out_0_839;
wire    [15:0]  conv_out_0_840, conv_out_0_841, conv_out_0_842, conv_out_0_843, conv_out_0_844, conv_out_0_845, conv_out_0_846, conv_out_0_847, conv_out_0_848, conv_out_0_849;
wire    [15:0]  conv_out_0_850, conv_out_0_851, conv_out_0_852, conv_out_0_853, conv_out_0_854, conv_out_0_855, conv_out_0_856, conv_out_0_857, conv_out_0_858, conv_out_0_859;
wire    [15:0]  conv_out_0_860, conv_out_0_861, conv_out_0_862, conv_out_0_863, conv_out_0_864, conv_out_0_865, conv_out_0_866, conv_out_0_867, conv_out_0_868, conv_out_0_869;
wire    [15:0]  conv_out_0_870, conv_out_0_871, conv_out_0_872, conv_out_0_873, conv_out_0_874, conv_out_0_875, conv_out_0_876, conv_out_0_877, conv_out_0_878, conv_out_0_879;
wire    [15:0]  conv_out_0_880, conv_out_0_881, conv_out_0_882, conv_out_0_883, conv_out_0_884, conv_out_0_885, conv_out_0_886, conv_out_0_887, conv_out_0_888, conv_out_0_889;
wire    [15:0]  conv_out_0_890, conv_out_0_891, conv_out_0_892, conv_out_0_893, conv_out_0_894, conv_out_0_895, conv_out_0_896, conv_out_0_897, conv_out_0_898, conv_out_0_899;

    
    wire    [35:0]  filter;

//    reg [15:0]  result  [899:0];

     assign  image_0_0[71:64]   = Image[0];
    assign  image_0_0[63:56]   = Image[1];
    assign  image_0_0[55:48]   = Image[2];
    assign  image_0_0[47:40]   = Image[32];
    assign  image_0_0[39:32]   = Image[33];
    assign  image_0_0[31:24]   = Image[34];
    assign  image_0_0[23:16]   = Image[64];
    assign  image_0_0[15:8]    = Image[65];
    assign  image_0_0[7:0]     = Image[66];

    assign  image_0_1[71:64]   = Image[1];
    assign  image_0_1[63:56]   = Image[2];
    assign  image_0_1[55:48]   = Image[3];
    assign  image_0_1[47:40]   = Image[33];
    assign  image_0_1[39:32]   = Image[34];
    assign  image_0_1[31:24]   = Image[35];
    assign  image_0_1[23:16]   = Image[65];
    assign  image_0_1[15:8]    = Image[66];
    assign  image_0_1[7:0]     = Image[67];

    assign  image_0_2[71:64]   = Image[2];
    assign  image_0_2[63:56]   = Image[3];
    assign  image_0_2[55:48]   = Image[4];
    assign  image_0_2[47:40]   = Image[34];
    assign  image_0_2[39:32]   = Image[35];
    assign  image_0_2[31:24]   = Image[36];
    assign  image_0_2[23:16]   = Image[66];
    assign  image_0_2[15:8]    = Image[67];
    assign  image_0_2[7:0]     = Image[68];

    assign  image_0_3[71:64]   = Image[3];
    assign  image_0_3[63:56]   = Image[4];
    assign  image_0_3[55:48]   = Image[5];
    assign  image_0_3[47:40]   = Image[35];
    assign  image_0_3[39:32]   = Image[36];
    assign  image_0_3[31:24]   = Image[37];
    assign  image_0_3[23:16]   = Image[67];
    assign  image_0_3[15:8]    = Image[68];
    assign  image_0_3[7:0]     = Image[69];

    assign  image_0_4[71:64]   = Image[4];
    assign  image_0_4[63:56]   = Image[5];
    assign  image_0_4[55:48]   = Image[6];
    assign  image_0_4[47:40]   = Image[36];
    assign  image_0_4[39:32]   = Image[37];
    assign  image_0_4[31:24]   = Image[38];
    assign  image_0_4[23:16]   = Image[68];
    assign  image_0_4[15:8]    = Image[69];
    assign  image_0_4[7:0]     = Image[70];

    assign  image_0_5[71:64]   = Image[5];
    assign  image_0_5[63:56]   = Image[6];
    assign  image_0_5[55:48]   = Image[7];
    assign  image_0_5[47:40]   = Image[37];
    assign  image_0_5[39:32]   = Image[38];
    assign  image_0_5[31:24]   = Image[39];
    assign  image_0_5[23:16]   = Image[69];
    assign  image_0_5[15:8]    = Image[70];
    assign  image_0_5[7:0]     = Image[71];

    assign  image_0_6[71:64]   = Image[6];
    assign  image_0_6[63:56]   = Image[7];
    assign  image_0_6[55:48]   = Image[8];
    assign  image_0_6[47:40]   = Image[38];
    assign  image_0_6[39:32]   = Image[39];
    assign  image_0_6[31:24]   = Image[40];
    assign  image_0_6[23:16]   = Image[70];
    assign  image_0_6[15:8]    = Image[71];
    assign  image_0_6[7:0]     = Image[72];

    assign  image_0_7[71:64]   = Image[7];
    assign  image_0_7[63:56]   = Image[8];
    assign  image_0_7[55:48]   = Image[9];
    assign  image_0_7[47:40]   = Image[39];
    assign  image_0_7[39:32]   = Image[40];
    assign  image_0_7[31:24]   = Image[41];
    assign  image_0_7[23:16]   = Image[71];
    assign  image_0_7[15:8]    = Image[72];
    assign  image_0_7[7:0]     = Image[73];

    assign  image_0_8[71:64]   = Image[8];
    assign  image_0_8[63:56]   = Image[9];
    assign  image_0_8[55:48]   = Image[10];
    assign  image_0_8[47:40]   = Image[40];
    assign  image_0_8[39:32]   = Image[41];
    assign  image_0_8[31:24]   = Image[42];
    assign  image_0_8[23:16]   = Image[72];
    assign  image_0_8[15:8]    = Image[73];
    assign  image_0_8[7:0]     = Image[74];

    assign  image_0_9[71:64]   = Image[9];
    assign  image_0_9[63:56]   = Image[10];
    assign  image_0_9[55:48]   = Image[11];
    assign  image_0_9[47:40]   = Image[41];
    assign  image_0_9[39:32]   = Image[42];
    assign  image_0_9[31:24]   = Image[43];
    assign  image_0_9[23:16]   = Image[73];
    assign  image_0_9[15:8]    = Image[74];
    assign  image_0_9[7:0]     = Image[75];

    assign  image_0_10[71:64]   = Image[10];
    assign  image_0_10[63:56]   = Image[11];
    assign  image_0_10[55:48]   = Image[12];
    assign  image_0_10[47:40]   = Image[42];
    assign  image_0_10[39:32]   = Image[43];
    assign  image_0_10[31:24]   = Image[44];
    assign  image_0_10[23:16]   = Image[74];
    assign  image_0_10[15:8]    = Image[75];
    assign  image_0_10[7:0]     = Image[76];

    assign  image_0_11[71:64]   = Image[11];
    assign  image_0_11[63:56]   = Image[12];
    assign  image_0_11[55:48]   = Image[13];
    assign  image_0_11[47:40]   = Image[43];
    assign  image_0_11[39:32]   = Image[44];
    assign  image_0_11[31:24]   = Image[45];
    assign  image_0_11[23:16]   = Image[75];
    assign  image_0_11[15:8]    = Image[76];
    assign  image_0_11[7:0]     = Image[77];

    assign  image_0_12[71:64]   = Image[12];
    assign  image_0_12[63:56]   = Image[13];
    assign  image_0_12[55:48]   = Image[14];
    assign  image_0_12[47:40]   = Image[44];
    assign  image_0_12[39:32]   = Image[45];
    assign  image_0_12[31:24]   = Image[46];
    assign  image_0_12[23:16]   = Image[76];
    assign  image_0_12[15:8]    = Image[77];
    assign  image_0_12[7:0]     = Image[78];

    assign  image_0_13[71:64]   = Image[13];
    assign  image_0_13[63:56]   = Image[14];
    assign  image_0_13[55:48]   = Image[15];
    assign  image_0_13[47:40]   = Image[45];
    assign  image_0_13[39:32]   = Image[46];
    assign  image_0_13[31:24]   = Image[47];
    assign  image_0_13[23:16]   = Image[77];
    assign  image_0_13[15:8]    = Image[78];
    assign  image_0_13[7:0]     = Image[79];

    assign  image_0_14[71:64]   = Image[14];
    assign  image_0_14[63:56]   = Image[15];
    assign  image_0_14[55:48]   = Image[16];
    assign  image_0_14[47:40]   = Image[46];
    assign  image_0_14[39:32]   = Image[47];
    assign  image_0_14[31:24]   = Image[48];
    assign  image_0_14[23:16]   = Image[78];
    assign  image_0_14[15:8]    = Image[79];
    assign  image_0_14[7:0]     = Image[80];

    assign  image_0_15[71:64]   = Image[15];
    assign  image_0_15[63:56]   = Image[16];
    assign  image_0_15[55:48]   = Image[17];
    assign  image_0_15[47:40]   = Image[47];
    assign  image_0_15[39:32]   = Image[48];
    assign  image_0_15[31:24]   = Image[49];
    assign  image_0_15[23:16]   = Image[79];
    assign  image_0_15[15:8]    = Image[80];
    assign  image_0_15[7:0]     = Image[81];

    assign  image_0_16[71:64]   = Image[16];
    assign  image_0_16[63:56]   = Image[17];
    assign  image_0_16[55:48]   = Image[18];
    assign  image_0_16[47:40]   = Image[48];
    assign  image_0_16[39:32]   = Image[49];
    assign  image_0_16[31:24]   = Image[50];
    assign  image_0_16[23:16]   = Image[80];
    assign  image_0_16[15:8]    = Image[81];
    assign  image_0_16[7:0]     = Image[82];

    assign  image_0_17[71:64]   = Image[17];
    assign  image_0_17[63:56]   = Image[18];
    assign  image_0_17[55:48]   = Image[19];
    assign  image_0_17[47:40]   = Image[49];
    assign  image_0_17[39:32]   = Image[50];
    assign  image_0_17[31:24]   = Image[51];
    assign  image_0_17[23:16]   = Image[81];
    assign  image_0_17[15:8]    = Image[82];
    assign  image_0_17[7:0]     = Image[83];

    assign  image_0_18[71:64]   = Image[18];
    assign  image_0_18[63:56]   = Image[19];
    assign  image_0_18[55:48]   = Image[20];
    assign  image_0_18[47:40]   = Image[50];
    assign  image_0_18[39:32]   = Image[51];
    assign  image_0_18[31:24]   = Image[52];
    assign  image_0_18[23:16]   = Image[82];
    assign  image_0_18[15:8]    = Image[83];
    assign  image_0_18[7:0]     = Image[84];

    assign  image_0_19[71:64]   = Image[19];
    assign  image_0_19[63:56]   = Image[20];
    assign  image_0_19[55:48]   = Image[21];
    assign  image_0_19[47:40]   = Image[51];
    assign  image_0_19[39:32]   = Image[52];
    assign  image_0_19[31:24]   = Image[53];
    assign  image_0_19[23:16]   = Image[83];
    assign  image_0_19[15:8]    = Image[84];
    assign  image_0_19[7:0]     = Image[85];

    assign  image_0_20[71:64]   = Image[20];
    assign  image_0_20[63:56]   = Image[21];
    assign  image_0_20[55:48]   = Image[22];
    assign  image_0_20[47:40]   = Image[52];
    assign  image_0_20[39:32]   = Image[53];
    assign  image_0_20[31:24]   = Image[54];
    assign  image_0_20[23:16]   = Image[84];
    assign  image_0_20[15:8]    = Image[85];
    assign  image_0_20[7:0]     = Image[86];

    assign  image_0_21[71:64]   = Image[21];
    assign  image_0_21[63:56]   = Image[22];
    assign  image_0_21[55:48]   = Image[23];
    assign  image_0_21[47:40]   = Image[53];
    assign  image_0_21[39:32]   = Image[54];
    assign  image_0_21[31:24]   = Image[55];
    assign  image_0_21[23:16]   = Image[85];
    assign  image_0_21[15:8]    = Image[86];
    assign  image_0_21[7:0]     = Image[87];

    assign  image_0_22[71:64]   = Image[22];
    assign  image_0_22[63:56]   = Image[23];
    assign  image_0_22[55:48]   = Image[24];
    assign  image_0_22[47:40]   = Image[54];
    assign  image_0_22[39:32]   = Image[55];
    assign  image_0_22[31:24]   = Image[56];
    assign  image_0_22[23:16]   = Image[86];
    assign  image_0_22[15:8]    = Image[87];
    assign  image_0_22[7:0]     = Image[88];

    assign  image_0_23[71:64]   = Image[23];
    assign  image_0_23[63:56]   = Image[24];
    assign  image_0_23[55:48]   = Image[25];
    assign  image_0_23[47:40]   = Image[55];
    assign  image_0_23[39:32]   = Image[56];
    assign  image_0_23[31:24]   = Image[57];
    assign  image_0_23[23:16]   = Image[87];
    assign  image_0_23[15:8]    = Image[88];
    assign  image_0_23[7:0]     = Image[89];

    assign  image_0_24[71:64]   = Image[24];
    assign  image_0_24[63:56]   = Image[25];
    assign  image_0_24[55:48]   = Image[26];
    assign  image_0_24[47:40]   = Image[56];
    assign  image_0_24[39:32]   = Image[57];
    assign  image_0_24[31:24]   = Image[58];
    assign  image_0_24[23:16]   = Image[88];
    assign  image_0_24[15:8]    = Image[89];
    assign  image_0_24[7:0]     = Image[90];

    assign  image_0_25[71:64]   = Image[25];
    assign  image_0_25[63:56]   = Image[26];
    assign  image_0_25[55:48]   = Image[27];
    assign  image_0_25[47:40]   = Image[57];
    assign  image_0_25[39:32]   = Image[58];
    assign  image_0_25[31:24]   = Image[59];
    assign  image_0_25[23:16]   = Image[89];
    assign  image_0_25[15:8]    = Image[90];
    assign  image_0_25[7:0]     = Image[91];

    assign  image_0_26[71:64]   = Image[26];
    assign  image_0_26[63:56]   = Image[27];
    assign  image_0_26[55:48]   = Image[28];
    assign  image_0_26[47:40]   = Image[58];
    assign  image_0_26[39:32]   = Image[59];
    assign  image_0_26[31:24]   = Image[60];
    assign  image_0_26[23:16]   = Image[90];
    assign  image_0_26[15:8]    = Image[91];
    assign  image_0_26[7:0]     = Image[92];

    assign  image_0_27[71:64]   = Image[27];
    assign  image_0_27[63:56]   = Image[28];
    assign  image_0_27[55:48]   = Image[29];
    assign  image_0_27[47:40]   = Image[59];
    assign  image_0_27[39:32]   = Image[60];
    assign  image_0_27[31:24]   = Image[61];
    assign  image_0_27[23:16]   = Image[91];
    assign  image_0_27[15:8]    = Image[92];
    assign  image_0_27[7:0]     = Image[93];

    assign  image_0_28[71:64]   = Image[28];
    assign  image_0_28[63:56]   = Image[29];
    assign  image_0_28[55:48]   = Image[30];
    assign  image_0_28[47:40]   = Image[60];
    assign  image_0_28[39:32]   = Image[61];
    assign  image_0_28[31:24]   = Image[62];
    assign  image_0_28[23:16]   = Image[92];
    assign  image_0_28[15:8]    = Image[93];
    assign  image_0_28[7:0]     = Image[94];

    assign  image_0_29[71:64]   = Image[29];
    assign  image_0_29[63:56]   = Image[30];
    assign  image_0_29[55:48]   = Image[31];
    assign  image_0_29[47:40]   = Image[61];
    assign  image_0_29[39:32]   = Image[62];
    assign  image_0_29[31:24]   = Image[63];
    assign  image_0_29[23:16]   = Image[93];
    assign  image_0_29[15:8]    = Image[94];
    assign  image_0_29[7:0]     = Image[95];

    assign  image_0_30[71:64]   = Image[32];
    assign  image_0_30[63:56]   = Image[33];
    assign  image_0_30[55:48]   = Image[34];
    assign  image_0_30[47:40]   = Image[64];
    assign  image_0_30[39:32]   = Image[65];
    assign  image_0_30[31:24]   = Image[66];
    assign  image_0_30[23:16]   = Image[96];
    assign  image_0_30[15:8]    = Image[97];
    assign  image_0_30[7:0]     = Image[98];

    assign  image_0_31[71:64]   = Image[33];
    assign  image_0_31[63:56]   = Image[34];
    assign  image_0_31[55:48]   = Image[35];
    assign  image_0_31[47:40]   = Image[65];
    assign  image_0_31[39:32]   = Image[66];
    assign  image_0_31[31:24]   = Image[67];
    assign  image_0_31[23:16]   = Image[97];
    assign  image_0_31[15:8]    = Image[98];
    assign  image_0_31[7:0]     = Image[99];

    assign  image_0_32[71:64]   = Image[34];
    assign  image_0_32[63:56]   = Image[35];
    assign  image_0_32[55:48]   = Image[36];
    assign  image_0_32[47:40]   = Image[66];
    assign  image_0_32[39:32]   = Image[67];
    assign  image_0_32[31:24]   = Image[68];
    assign  image_0_32[23:16]   = Image[98];
    assign  image_0_32[15:8]    = Image[99];
    assign  image_0_32[7:0]     = Image[100];

    assign  image_0_33[71:64]   = Image[35];
    assign  image_0_33[63:56]   = Image[36];
    assign  image_0_33[55:48]   = Image[37];
    assign  image_0_33[47:40]   = Image[67];
    assign  image_0_33[39:32]   = Image[68];
    assign  image_0_33[31:24]   = Image[69];
    assign  image_0_33[23:16]   = Image[99];
    assign  image_0_33[15:8]    = Image[100];
    assign  image_0_33[7:0]     = Image[101];

    assign  image_0_34[71:64]   = Image[36];
    assign  image_0_34[63:56]   = Image[37];
    assign  image_0_34[55:48]   = Image[38];
    assign  image_0_34[47:40]   = Image[68];
    assign  image_0_34[39:32]   = Image[69];
    assign  image_0_34[31:24]   = Image[70];
    assign  image_0_34[23:16]   = Image[100];
    assign  image_0_34[15:8]    = Image[101];
    assign  image_0_34[7:0]     = Image[102];

    assign  image_0_35[71:64]   = Image[37];
    assign  image_0_35[63:56]   = Image[38];
    assign  image_0_35[55:48]   = Image[39];
    assign  image_0_35[47:40]   = Image[69];
    assign  image_0_35[39:32]   = Image[70];
    assign  image_0_35[31:24]   = Image[71];
    assign  image_0_35[23:16]   = Image[101];
    assign  image_0_35[15:8]    = Image[102];
    assign  image_0_35[7:0]     = Image[103];

    assign  image_0_36[71:64]   = Image[38];
    assign  image_0_36[63:56]   = Image[39];
    assign  image_0_36[55:48]   = Image[40];
    assign  image_0_36[47:40]   = Image[70];
    assign  image_0_36[39:32]   = Image[71];
    assign  image_0_36[31:24]   = Image[72];
    assign  image_0_36[23:16]   = Image[102];
    assign  image_0_36[15:8]    = Image[103];
    assign  image_0_36[7:0]     = Image[104];

    assign  image_0_37[71:64]   = Image[39];
    assign  image_0_37[63:56]   = Image[40];
    assign  image_0_37[55:48]   = Image[41];
    assign  image_0_37[47:40]   = Image[71];
    assign  image_0_37[39:32]   = Image[72];
    assign  image_0_37[31:24]   = Image[73];
    assign  image_0_37[23:16]   = Image[103];
    assign  image_0_37[15:8]    = Image[104];
    assign  image_0_37[7:0]     = Image[105];

    assign  image_0_38[71:64]   = Image[40];
    assign  image_0_38[63:56]   = Image[41];
    assign  image_0_38[55:48]   = Image[42];
    assign  image_0_38[47:40]   = Image[72];
    assign  image_0_38[39:32]   = Image[73];
    assign  image_0_38[31:24]   = Image[74];
    assign  image_0_38[23:16]   = Image[104];
    assign  image_0_38[15:8]    = Image[105];
    assign  image_0_38[7:0]     = Image[106];

    assign  image_0_39[71:64]   = Image[41];
    assign  image_0_39[63:56]   = Image[42];
    assign  image_0_39[55:48]   = Image[43];
    assign  image_0_39[47:40]   = Image[73];
    assign  image_0_39[39:32]   = Image[74];
    assign  image_0_39[31:24]   = Image[75];
    assign  image_0_39[23:16]   = Image[105];
    assign  image_0_39[15:8]    = Image[106];
    assign  image_0_39[7:0]     = Image[107];

    assign  image_0_40[71:64]   = Image[42];
    assign  image_0_40[63:56]   = Image[43];
    assign  image_0_40[55:48]   = Image[44];
    assign  image_0_40[47:40]   = Image[74];
    assign  image_0_40[39:32]   = Image[75];
    assign  image_0_40[31:24]   = Image[76];
    assign  image_0_40[23:16]   = Image[106];
    assign  image_0_40[15:8]    = Image[107];
    assign  image_0_40[7:0]     = Image[108];

    assign  image_0_41[71:64]   = Image[43];
    assign  image_0_41[63:56]   = Image[44];
    assign  image_0_41[55:48]   = Image[45];
    assign  image_0_41[47:40]   = Image[75];
    assign  image_0_41[39:32]   = Image[76];
    assign  image_0_41[31:24]   = Image[77];
    assign  image_0_41[23:16]   = Image[107];
    assign  image_0_41[15:8]    = Image[108];
    assign  image_0_41[7:0]     = Image[109];

    assign  image_0_42[71:64]   = Image[44];
    assign  image_0_42[63:56]   = Image[45];
    assign  image_0_42[55:48]   = Image[46];
    assign  image_0_42[47:40]   = Image[76];
    assign  image_0_42[39:32]   = Image[77];
    assign  image_0_42[31:24]   = Image[78];
    assign  image_0_42[23:16]   = Image[108];
    assign  image_0_42[15:8]    = Image[109];
    assign  image_0_42[7:0]     = Image[110];

    assign  image_0_43[71:64]   = Image[45];
    assign  image_0_43[63:56]   = Image[46];
    assign  image_0_43[55:48]   = Image[47];
    assign  image_0_43[47:40]   = Image[77];
    assign  image_0_43[39:32]   = Image[78];
    assign  image_0_43[31:24]   = Image[79];
    assign  image_0_43[23:16]   = Image[109];
    assign  image_0_43[15:8]    = Image[110];
    assign  image_0_43[7:0]     = Image[111];

    assign  image_0_44[71:64]   = Image[46];
    assign  image_0_44[63:56]   = Image[47];
    assign  image_0_44[55:48]   = Image[48];
    assign  image_0_44[47:40]   = Image[78];
    assign  image_0_44[39:32]   = Image[79];
    assign  image_0_44[31:24]   = Image[80];
    assign  image_0_44[23:16]   = Image[110];
    assign  image_0_44[15:8]    = Image[111];
    assign  image_0_44[7:0]     = Image[112];

    assign  image_0_45[71:64]   = Image[47];
    assign  image_0_45[63:56]   = Image[48];
    assign  image_0_45[55:48]   = Image[49];
    assign  image_0_45[47:40]   = Image[79];
    assign  image_0_45[39:32]   = Image[80];
    assign  image_0_45[31:24]   = Image[81];
    assign  image_0_45[23:16]   = Image[111];
    assign  image_0_45[15:8]    = Image[112];
    assign  image_0_45[7:0]     = Image[113];

    assign  image_0_46[71:64]   = Image[48];
    assign  image_0_46[63:56]   = Image[49];
    assign  image_0_46[55:48]   = Image[50];
    assign  image_0_46[47:40]   = Image[80];
    assign  image_0_46[39:32]   = Image[81];
    assign  image_0_46[31:24]   = Image[82];
    assign  image_0_46[23:16]   = Image[112];
    assign  image_0_46[15:8]    = Image[113];
    assign  image_0_46[7:0]     = Image[114];

    assign  image_0_47[71:64]   = Image[49];
    assign  image_0_47[63:56]   = Image[50];
    assign  image_0_47[55:48]   = Image[51];
    assign  image_0_47[47:40]   = Image[81];
    assign  image_0_47[39:32]   = Image[82];
    assign  image_0_47[31:24]   = Image[83];
    assign  image_0_47[23:16]   = Image[113];
    assign  image_0_47[15:8]    = Image[114];
    assign  image_0_47[7:0]     = Image[115];

    assign  image_0_48[71:64]   = Image[50];
    assign  image_0_48[63:56]   = Image[51];
    assign  image_0_48[55:48]   = Image[52];
    assign  image_0_48[47:40]   = Image[82];
    assign  image_0_48[39:32]   = Image[83];
    assign  image_0_48[31:24]   = Image[84];
    assign  image_0_48[23:16]   = Image[114];
    assign  image_0_48[15:8]    = Image[115];
    assign  image_0_48[7:0]     = Image[116];

    assign  image_0_49[71:64]   = Image[51];
    assign  image_0_49[63:56]   = Image[52];
    assign  image_0_49[55:48]   = Image[53];
    assign  image_0_49[47:40]   = Image[83];
    assign  image_0_49[39:32]   = Image[84];
    assign  image_0_49[31:24]   = Image[85];
    assign  image_0_49[23:16]   = Image[115];
    assign  image_0_49[15:8]    = Image[116];
    assign  image_0_49[7:0]     = Image[117];

    assign  image_0_50[71:64]   = Image[52];
    assign  image_0_50[63:56]   = Image[53];
    assign  image_0_50[55:48]   = Image[54];
    assign  image_0_50[47:40]   = Image[84];
    assign  image_0_50[39:32]   = Image[85];
    assign  image_0_50[31:24]   = Image[86];
    assign  image_0_50[23:16]   = Image[116];
    assign  image_0_50[15:8]    = Image[117];
    assign  image_0_50[7:0]     = Image[118];

    assign  image_0_51[71:64]   = Image[53];
    assign  image_0_51[63:56]   = Image[54];
    assign  image_0_51[55:48]   = Image[55];
    assign  image_0_51[47:40]   = Image[85];
    assign  image_0_51[39:32]   = Image[86];
    assign  image_0_51[31:24]   = Image[87];
    assign  image_0_51[23:16]   = Image[117];
    assign  image_0_51[15:8]    = Image[118];
    assign  image_0_51[7:0]     = Image[119];

    assign  image_0_52[71:64]   = Image[54];
    assign  image_0_52[63:56]   = Image[55];
    assign  image_0_52[55:48]   = Image[56];
    assign  image_0_52[47:40]   = Image[86];
    assign  image_0_52[39:32]   = Image[87];
    assign  image_0_52[31:24]   = Image[88];
    assign  image_0_52[23:16]   = Image[118];
    assign  image_0_52[15:8]    = Image[119];
    assign  image_0_52[7:0]     = Image[120];

    assign  image_0_53[71:64]   = Image[55];
    assign  image_0_53[63:56]   = Image[56];
    assign  image_0_53[55:48]   = Image[57];
    assign  image_0_53[47:40]   = Image[87];
    assign  image_0_53[39:32]   = Image[88];
    assign  image_0_53[31:24]   = Image[89];
    assign  image_0_53[23:16]   = Image[119];
    assign  image_0_53[15:8]    = Image[120];
    assign  image_0_53[7:0]     = Image[121];

    assign  image_0_54[71:64]   = Image[56];
    assign  image_0_54[63:56]   = Image[57];
    assign  image_0_54[55:48]   = Image[58];
    assign  image_0_54[47:40]   = Image[88];
    assign  image_0_54[39:32]   = Image[89];
    assign  image_0_54[31:24]   = Image[90];
    assign  image_0_54[23:16]   = Image[120];
    assign  image_0_54[15:8]    = Image[121];
    assign  image_0_54[7:0]     = Image[122];

    assign  image_0_55[71:64]   = Image[57];
    assign  image_0_55[63:56]   = Image[58];
    assign  image_0_55[55:48]   = Image[59];
    assign  image_0_55[47:40]   = Image[89];
    assign  image_0_55[39:32]   = Image[90];
    assign  image_0_55[31:24]   = Image[91];
    assign  image_0_55[23:16]   = Image[121];
    assign  image_0_55[15:8]    = Image[122];
    assign  image_0_55[7:0]     = Image[123];

    assign  image_0_56[71:64]   = Image[58];
    assign  image_0_56[63:56]   = Image[59];
    assign  image_0_56[55:48]   = Image[60];
    assign  image_0_56[47:40]   = Image[90];
    assign  image_0_56[39:32]   = Image[91];
    assign  image_0_56[31:24]   = Image[92];
    assign  image_0_56[23:16]   = Image[122];
    assign  image_0_56[15:8]    = Image[123];
    assign  image_0_56[7:0]     = Image[124];

    assign  image_0_57[71:64]   = Image[59];
    assign  image_0_57[63:56]   = Image[60];
    assign  image_0_57[55:48]   = Image[61];
    assign  image_0_57[47:40]   = Image[91];
    assign  image_0_57[39:32]   = Image[92];
    assign  image_0_57[31:24]   = Image[93];
    assign  image_0_57[23:16]   = Image[123];
    assign  image_0_57[15:8]    = Image[124];
    assign  image_0_57[7:0]     = Image[125];

    assign  image_0_58[71:64]   = Image[60];
    assign  image_0_58[63:56]   = Image[61];
    assign  image_0_58[55:48]   = Image[62];
    assign  image_0_58[47:40]   = Image[92];
    assign  image_0_58[39:32]   = Image[93];
    assign  image_0_58[31:24]   = Image[94];
    assign  image_0_58[23:16]   = Image[124];
    assign  image_0_58[15:8]    = Image[125];
    assign  image_0_58[7:0]     = Image[126];

    assign  image_0_59[71:64]   = Image[61];
    assign  image_0_59[63:56]   = Image[62];
    assign  image_0_59[55:48]   = Image[63];
    assign  image_0_59[47:40]   = Image[93];
    assign  image_0_59[39:32]   = Image[94];
    assign  image_0_59[31:24]   = Image[95];
    assign  image_0_59[23:16]   = Image[125];
    assign  image_0_59[15:8]    = Image[126];
    assign  image_0_59[7:0]     = Image[127];

    assign  image_0_60[71:64]   = Image[64];
    assign  image_0_60[63:56]   = Image[65];
    assign  image_0_60[55:48]   = Image[66];
    assign  image_0_60[47:40]   = Image[96];
    assign  image_0_60[39:32]   = Image[97];
    assign  image_0_60[31:24]   = Image[98];
    assign  image_0_60[23:16]   = Image[128];
    assign  image_0_60[15:8]    = Image[129];
    assign  image_0_60[7:0]     = Image[130];

    assign  image_0_61[71:64]   = Image[65];
    assign  image_0_61[63:56]   = Image[66];
    assign  image_0_61[55:48]   = Image[67];
    assign  image_0_61[47:40]   = Image[97];
    assign  image_0_61[39:32]   = Image[98];
    assign  image_0_61[31:24]   = Image[99];
    assign  image_0_61[23:16]   = Image[129];
    assign  image_0_61[15:8]    = Image[130];
    assign  image_0_61[7:0]     = Image[131];

    assign  image_0_62[71:64]   = Image[66];
    assign  image_0_62[63:56]   = Image[67];
    assign  image_0_62[55:48]   = Image[68];
    assign  image_0_62[47:40]   = Image[98];
    assign  image_0_62[39:32]   = Image[99];
    assign  image_0_62[31:24]   = Image[100];
    assign  image_0_62[23:16]   = Image[130];
    assign  image_0_62[15:8]    = Image[131];
    assign  image_0_62[7:0]     = Image[132];

    assign  image_0_63[71:64]   = Image[67];
    assign  image_0_63[63:56]   = Image[68];
    assign  image_0_63[55:48]   = Image[69];
    assign  image_0_63[47:40]   = Image[99];
    assign  image_0_63[39:32]   = Image[100];
    assign  image_0_63[31:24]   = Image[101];
    assign  image_0_63[23:16]   = Image[131];
    assign  image_0_63[15:8]    = Image[132];
    assign  image_0_63[7:0]     = Image[133];

    assign  image_0_64[71:64]   = Image[68];
    assign  image_0_64[63:56]   = Image[69];
    assign  image_0_64[55:48]   = Image[70];
    assign  image_0_64[47:40]   = Image[100];
    assign  image_0_64[39:32]   = Image[101];
    assign  image_0_64[31:24]   = Image[102];
    assign  image_0_64[23:16]   = Image[132];
    assign  image_0_64[15:8]    = Image[133];
    assign  image_0_64[7:0]     = Image[134];

    assign  image_0_65[71:64]   = Image[69];
    assign  image_0_65[63:56]   = Image[70];
    assign  image_0_65[55:48]   = Image[71];
    assign  image_0_65[47:40]   = Image[101];
    assign  image_0_65[39:32]   = Image[102];
    assign  image_0_65[31:24]   = Image[103];
    assign  image_0_65[23:16]   = Image[133];
    assign  image_0_65[15:8]    = Image[134];
    assign  image_0_65[7:0]     = Image[135];

    assign  image_0_66[71:64]   = Image[70];
    assign  image_0_66[63:56]   = Image[71];
    assign  image_0_66[55:48]   = Image[72];
    assign  image_0_66[47:40]   = Image[102];
    assign  image_0_66[39:32]   = Image[103];
    assign  image_0_66[31:24]   = Image[104];
    assign  image_0_66[23:16]   = Image[134];
    assign  image_0_66[15:8]    = Image[135];
    assign  image_0_66[7:0]     = Image[136];

    assign  image_0_67[71:64]   = Image[71];
    assign  image_0_67[63:56]   = Image[72];
    assign  image_0_67[55:48]   = Image[73];
    assign  image_0_67[47:40]   = Image[103];
    assign  image_0_67[39:32]   = Image[104];
    assign  image_0_67[31:24]   = Image[105];
    assign  image_0_67[23:16]   = Image[135];
    assign  image_0_67[15:8]    = Image[136];
    assign  image_0_67[7:0]     = Image[137];

    assign  image_0_68[71:64]   = Image[72];
    assign  image_0_68[63:56]   = Image[73];
    assign  image_0_68[55:48]   = Image[74];
    assign  image_0_68[47:40]   = Image[104];
    assign  image_0_68[39:32]   = Image[105];
    assign  image_0_68[31:24]   = Image[106];
    assign  image_0_68[23:16]   = Image[136];
    assign  image_0_68[15:8]    = Image[137];
    assign  image_0_68[7:0]     = Image[138];

    assign  image_0_69[71:64]   = Image[73];
    assign  image_0_69[63:56]   = Image[74];
    assign  image_0_69[55:48]   = Image[75];
    assign  image_0_69[47:40]   = Image[105];
    assign  image_0_69[39:32]   = Image[106];
    assign  image_0_69[31:24]   = Image[107];
    assign  image_0_69[23:16]   = Image[137];
    assign  image_0_69[15:8]    = Image[138];
    assign  image_0_69[7:0]     = Image[139];

    assign  image_0_70[71:64]   = Image[74];
    assign  image_0_70[63:56]   = Image[75];
    assign  image_0_70[55:48]   = Image[76];
    assign  image_0_70[47:40]   = Image[106];
    assign  image_0_70[39:32]   = Image[107];
    assign  image_0_70[31:24]   = Image[108];
    assign  image_0_70[23:16]   = Image[138];
    assign  image_0_70[15:8]    = Image[139];
    assign  image_0_70[7:0]     = Image[140];

    assign  image_0_71[71:64]   = Image[75];
    assign  image_0_71[63:56]   = Image[76];
    assign  image_0_71[55:48]   = Image[77];
    assign  image_0_71[47:40]   = Image[107];
    assign  image_0_71[39:32]   = Image[108];
    assign  image_0_71[31:24]   = Image[109];
    assign  image_0_71[23:16]   = Image[139];
    assign  image_0_71[15:8]    = Image[140];
    assign  image_0_71[7:0]     = Image[141];

    assign  image_0_72[71:64]   = Image[76];
    assign  image_0_72[63:56]   = Image[77];
    assign  image_0_72[55:48]   = Image[78];
    assign  image_0_72[47:40]   = Image[108];
    assign  image_0_72[39:32]   = Image[109];
    assign  image_0_72[31:24]   = Image[110];
    assign  image_0_72[23:16]   = Image[140];
    assign  image_0_72[15:8]    = Image[141];
    assign  image_0_72[7:0]     = Image[142];

    assign  image_0_73[71:64]   = Image[77];
    assign  image_0_73[63:56]   = Image[78];
    assign  image_0_73[55:48]   = Image[79];
    assign  image_0_73[47:40]   = Image[109];
    assign  image_0_73[39:32]   = Image[110];
    assign  image_0_73[31:24]   = Image[111];
    assign  image_0_73[23:16]   = Image[141];
    assign  image_0_73[15:8]    = Image[142];
    assign  image_0_73[7:0]     = Image[143];

    assign  image_0_74[71:64]   = Image[78];
    assign  image_0_74[63:56]   = Image[79];
    assign  image_0_74[55:48]   = Image[80];
    assign  image_0_74[47:40]   = Image[110];
    assign  image_0_74[39:32]   = Image[111];
    assign  image_0_74[31:24]   = Image[112];
    assign  image_0_74[23:16]   = Image[142];
    assign  image_0_74[15:8]    = Image[143];
    assign  image_0_74[7:0]     = Image[144];

    assign  image_0_75[71:64]   = Image[79];
    assign  image_0_75[63:56]   = Image[80];
    assign  image_0_75[55:48]   = Image[81];
    assign  image_0_75[47:40]   = Image[111];
    assign  image_0_75[39:32]   = Image[112];
    assign  image_0_75[31:24]   = Image[113];
    assign  image_0_75[23:16]   = Image[143];
    assign  image_0_75[15:8]    = Image[144];
    assign  image_0_75[7:0]     = Image[145];

    assign  image_0_76[71:64]   = Image[80];
    assign  image_0_76[63:56]   = Image[81];
    assign  image_0_76[55:48]   = Image[82];
    assign  image_0_76[47:40]   = Image[112];
    assign  image_0_76[39:32]   = Image[113];
    assign  image_0_76[31:24]   = Image[114];
    assign  image_0_76[23:16]   = Image[144];
    assign  image_0_76[15:8]    = Image[145];
    assign  image_0_76[7:0]     = Image[146];

    assign  image_0_77[71:64]   = Image[81];
    assign  image_0_77[63:56]   = Image[82];
    assign  image_0_77[55:48]   = Image[83];
    assign  image_0_77[47:40]   = Image[113];
    assign  image_0_77[39:32]   = Image[114];
    assign  image_0_77[31:24]   = Image[115];
    assign  image_0_77[23:16]   = Image[145];
    assign  image_0_77[15:8]    = Image[146];
    assign  image_0_77[7:0]     = Image[147];

    assign  image_0_78[71:64]   = Image[82];
    assign  image_0_78[63:56]   = Image[83];
    assign  image_0_78[55:48]   = Image[84];
    assign  image_0_78[47:40]   = Image[114];
    assign  image_0_78[39:32]   = Image[115];
    assign  image_0_78[31:24]   = Image[116];
    assign  image_0_78[23:16]   = Image[146];
    assign  image_0_78[15:8]    = Image[147];
    assign  image_0_78[7:0]     = Image[148];

    assign  image_0_79[71:64]   = Image[83];
    assign  image_0_79[63:56]   = Image[84];
    assign  image_0_79[55:48]   = Image[85];
    assign  image_0_79[47:40]   = Image[115];
    assign  image_0_79[39:32]   = Image[116];
    assign  image_0_79[31:24]   = Image[117];
    assign  image_0_79[23:16]   = Image[147];
    assign  image_0_79[15:8]    = Image[148];
    assign  image_0_79[7:0]     = Image[149];

    assign  image_0_80[71:64]   = Image[84];
    assign  image_0_80[63:56]   = Image[85];
    assign  image_0_80[55:48]   = Image[86];
    assign  image_0_80[47:40]   = Image[116];
    assign  image_0_80[39:32]   = Image[117];
    assign  image_0_80[31:24]   = Image[118];
    assign  image_0_80[23:16]   = Image[148];
    assign  image_0_80[15:8]    = Image[149];
    assign  image_0_80[7:0]     = Image[150];

    assign  image_0_81[71:64]   = Image[85];
    assign  image_0_81[63:56]   = Image[86];
    assign  image_0_81[55:48]   = Image[87];
    assign  image_0_81[47:40]   = Image[117];
    assign  image_0_81[39:32]   = Image[118];
    assign  image_0_81[31:24]   = Image[119];
    assign  image_0_81[23:16]   = Image[149];
    assign  image_0_81[15:8]    = Image[150];
    assign  image_0_81[7:0]     = Image[151];

    assign  image_0_82[71:64]   = Image[86];
    assign  image_0_82[63:56]   = Image[87];
    assign  image_0_82[55:48]   = Image[88];
    assign  image_0_82[47:40]   = Image[118];
    assign  image_0_82[39:32]   = Image[119];
    assign  image_0_82[31:24]   = Image[120];
    assign  image_0_82[23:16]   = Image[150];
    assign  image_0_82[15:8]    = Image[151];
    assign  image_0_82[7:0]     = Image[152];

    assign  image_0_83[71:64]   = Image[87];
    assign  image_0_83[63:56]   = Image[88];
    assign  image_0_83[55:48]   = Image[89];
    assign  image_0_83[47:40]   = Image[119];
    assign  image_0_83[39:32]   = Image[120];
    assign  image_0_83[31:24]   = Image[121];
    assign  image_0_83[23:16]   = Image[151];
    assign  image_0_83[15:8]    = Image[152];
    assign  image_0_83[7:0]     = Image[153];

    assign  image_0_84[71:64]   = Image[88];
    assign  image_0_84[63:56]   = Image[89];
    assign  image_0_84[55:48]   = Image[90];
    assign  image_0_84[47:40]   = Image[120];
    assign  image_0_84[39:32]   = Image[121];
    assign  image_0_84[31:24]   = Image[122];
    assign  image_0_84[23:16]   = Image[152];
    assign  image_0_84[15:8]    = Image[153];
    assign  image_0_84[7:0]     = Image[154];

    assign  image_0_85[71:64]   = Image[89];
    assign  image_0_85[63:56]   = Image[90];
    assign  image_0_85[55:48]   = Image[91];
    assign  image_0_85[47:40]   = Image[121];
    assign  image_0_85[39:32]   = Image[122];
    assign  image_0_85[31:24]   = Image[123];
    assign  image_0_85[23:16]   = Image[153];
    assign  image_0_85[15:8]    = Image[154];
    assign  image_0_85[7:0]     = Image[155];

    assign  image_0_86[71:64]   = Image[90];
    assign  image_0_86[63:56]   = Image[91];
    assign  image_0_86[55:48]   = Image[92];
    assign  image_0_86[47:40]   = Image[122];
    assign  image_0_86[39:32]   = Image[123];
    assign  image_0_86[31:24]   = Image[124];
    assign  image_0_86[23:16]   = Image[154];
    assign  image_0_86[15:8]    = Image[155];
    assign  image_0_86[7:0]     = Image[156];

    assign  image_0_87[71:64]   = Image[91];
    assign  image_0_87[63:56]   = Image[92];
    assign  image_0_87[55:48]   = Image[93];
    assign  image_0_87[47:40]   = Image[123];
    assign  image_0_87[39:32]   = Image[124];
    assign  image_0_87[31:24]   = Image[125];
    assign  image_0_87[23:16]   = Image[155];
    assign  image_0_87[15:8]    = Image[156];
    assign  image_0_87[7:0]     = Image[157];

    assign  image_0_88[71:64]   = Image[92];
    assign  image_0_88[63:56]   = Image[93];
    assign  image_0_88[55:48]   = Image[94];
    assign  image_0_88[47:40]   = Image[124];
    assign  image_0_88[39:32]   = Image[125];
    assign  image_0_88[31:24]   = Image[126];
    assign  image_0_88[23:16]   = Image[156];
    assign  image_0_88[15:8]    = Image[157];
    assign  image_0_88[7:0]     = Image[158];

    assign  image_0_89[71:64]   = Image[93];
    assign  image_0_89[63:56]   = Image[94];
    assign  image_0_89[55:48]   = Image[95];
    assign  image_0_89[47:40]   = Image[125];
    assign  image_0_89[39:32]   = Image[126];
    assign  image_0_89[31:24]   = Image[127];
    assign  image_0_89[23:16]   = Image[157];
    assign  image_0_89[15:8]    = Image[158];
    assign  image_0_89[7:0]     = Image[159];

    assign  image_0_90[71:64]   = Image[96];
    assign  image_0_90[63:56]   = Image[97];
    assign  image_0_90[55:48]   = Image[98];
    assign  image_0_90[47:40]   = Image[128];
    assign  image_0_90[39:32]   = Image[129];
    assign  image_0_90[31:24]   = Image[130];
    assign  image_0_90[23:16]   = Image[160];
    assign  image_0_90[15:8]    = Image[161];
    assign  image_0_90[7:0]     = Image[162];

    assign  image_0_91[71:64]   = Image[97];
    assign  image_0_91[63:56]   = Image[98];
    assign  image_0_91[55:48]   = Image[99];
    assign  image_0_91[47:40]   = Image[129];
    assign  image_0_91[39:32]   = Image[130];
    assign  image_0_91[31:24]   = Image[131];
    assign  image_0_91[23:16]   = Image[161];
    assign  image_0_91[15:8]    = Image[162];
    assign  image_0_91[7:0]     = Image[163];

    assign  image_0_92[71:64]   = Image[98];
    assign  image_0_92[63:56]   = Image[99];
    assign  image_0_92[55:48]   = Image[100];
    assign  image_0_92[47:40]   = Image[130];
    assign  image_0_92[39:32]   = Image[131];
    assign  image_0_92[31:24]   = Image[132];
    assign  image_0_92[23:16]   = Image[162];
    assign  image_0_92[15:8]    = Image[163];
    assign  image_0_92[7:0]     = Image[164];

    assign  image_0_93[71:64]   = Image[99];
    assign  image_0_93[63:56]   = Image[100];
    assign  image_0_93[55:48]   = Image[101];
    assign  image_0_93[47:40]   = Image[131];
    assign  image_0_93[39:32]   = Image[132];
    assign  image_0_93[31:24]   = Image[133];
    assign  image_0_93[23:16]   = Image[163];
    assign  image_0_93[15:8]    = Image[164];
    assign  image_0_93[7:0]     = Image[165];

    assign  image_0_94[71:64]   = Image[100];
    assign  image_0_94[63:56]   = Image[101];
    assign  image_0_94[55:48]   = Image[102];
    assign  image_0_94[47:40]   = Image[132];
    assign  image_0_94[39:32]   = Image[133];
    assign  image_0_94[31:24]   = Image[134];
    assign  image_0_94[23:16]   = Image[164];
    assign  image_0_94[15:8]    = Image[165];
    assign  image_0_94[7:0]     = Image[166];

    assign  image_0_95[71:64]   = Image[101];
    assign  image_0_95[63:56]   = Image[102];
    assign  image_0_95[55:48]   = Image[103];
    assign  image_0_95[47:40]   = Image[133];
    assign  image_0_95[39:32]   = Image[134];
    assign  image_0_95[31:24]   = Image[135];
    assign  image_0_95[23:16]   = Image[165];
    assign  image_0_95[15:8]    = Image[166];
    assign  image_0_95[7:0]     = Image[167];

    assign  image_0_96[71:64]   = Image[102];
    assign  image_0_96[63:56]   = Image[103];
    assign  image_0_96[55:48]   = Image[104];
    assign  image_0_96[47:40]   = Image[134];
    assign  image_0_96[39:32]   = Image[135];
    assign  image_0_96[31:24]   = Image[136];
    assign  image_0_96[23:16]   = Image[166];
    assign  image_0_96[15:8]    = Image[167];
    assign  image_0_96[7:0]     = Image[168];

    assign  image_0_97[71:64]   = Image[103];
    assign  image_0_97[63:56]   = Image[104];
    assign  image_0_97[55:48]   = Image[105];
    assign  image_0_97[47:40]   = Image[135];
    assign  image_0_97[39:32]   = Image[136];
    assign  image_0_97[31:24]   = Image[137];
    assign  image_0_97[23:16]   = Image[167];
    assign  image_0_97[15:8]    = Image[168];
    assign  image_0_97[7:0]     = Image[169];

    assign  image_0_98[71:64]   = Image[104];
    assign  image_0_98[63:56]   = Image[105];
    assign  image_0_98[55:48]   = Image[106];
    assign  image_0_98[47:40]   = Image[136];
    assign  image_0_98[39:32]   = Image[137];
    assign  image_0_98[31:24]   = Image[138];
    assign  image_0_98[23:16]   = Image[168];
    assign  image_0_98[15:8]    = Image[169];
    assign  image_0_98[7:0]     = Image[170];

    assign  image_0_99[71:64]   = Image[105];
    assign  image_0_99[63:56]   = Image[106];
    assign  image_0_99[55:48]   = Image[107];
    assign  image_0_99[47:40]   = Image[137];
    assign  image_0_99[39:32]   = Image[138];
    assign  image_0_99[31:24]   = Image[139];
    assign  image_0_99[23:16]   = Image[169];
    assign  image_0_99[15:8]    = Image[170];
    assign  image_0_99[7:0]     = Image[171];

    assign  image_0_100[71:64]   = Image[106];
    assign  image_0_100[63:56]   = Image[107];
    assign  image_0_100[55:48]   = Image[108];
    assign  image_0_100[47:40]   = Image[138];
    assign  image_0_100[39:32]   = Image[139];
    assign  image_0_100[31:24]   = Image[140];
    assign  image_0_100[23:16]   = Image[170];
    assign  image_0_100[15:8]    = Image[171];
    assign  image_0_100[7:0]     = Image[172];

    assign  image_0_101[71:64]   = Image[107];
    assign  image_0_101[63:56]   = Image[108];
    assign  image_0_101[55:48]   = Image[109];
    assign  image_0_101[47:40]   = Image[139];
    assign  image_0_101[39:32]   = Image[140];
    assign  image_0_101[31:24]   = Image[141];
    assign  image_0_101[23:16]   = Image[171];
    assign  image_0_101[15:8]    = Image[172];
    assign  image_0_101[7:0]     = Image[173];

    assign  image_0_102[71:64]   = Image[108];
    assign  image_0_102[63:56]   = Image[109];
    assign  image_0_102[55:48]   = Image[110];
    assign  image_0_102[47:40]   = Image[140];
    assign  image_0_102[39:32]   = Image[141];
    assign  image_0_102[31:24]   = Image[142];
    assign  image_0_102[23:16]   = Image[172];
    assign  image_0_102[15:8]    = Image[173];
    assign  image_0_102[7:0]     = Image[174];

    assign  image_0_103[71:64]   = Image[109];
    assign  image_0_103[63:56]   = Image[110];
    assign  image_0_103[55:48]   = Image[111];
    assign  image_0_103[47:40]   = Image[141];
    assign  image_0_103[39:32]   = Image[142];
    assign  image_0_103[31:24]   = Image[143];
    assign  image_0_103[23:16]   = Image[173];
    assign  image_0_103[15:8]    = Image[174];
    assign  image_0_103[7:0]     = Image[175];

    assign  image_0_104[71:64]   = Image[110];
    assign  image_0_104[63:56]   = Image[111];
    assign  image_0_104[55:48]   = Image[112];
    assign  image_0_104[47:40]   = Image[142];
    assign  image_0_104[39:32]   = Image[143];
    assign  image_0_104[31:24]   = Image[144];
    assign  image_0_104[23:16]   = Image[174];
    assign  image_0_104[15:8]    = Image[175];
    assign  image_0_104[7:0]     = Image[176];

    assign  image_0_105[71:64]   = Image[111];
    assign  image_0_105[63:56]   = Image[112];
    assign  image_0_105[55:48]   = Image[113];
    assign  image_0_105[47:40]   = Image[143];
    assign  image_0_105[39:32]   = Image[144];
    assign  image_0_105[31:24]   = Image[145];
    assign  image_0_105[23:16]   = Image[175];
    assign  image_0_105[15:8]    = Image[176];
    assign  image_0_105[7:0]     = Image[177];

    assign  image_0_106[71:64]   = Image[112];
    assign  image_0_106[63:56]   = Image[113];
    assign  image_0_106[55:48]   = Image[114];
    assign  image_0_106[47:40]   = Image[144];
    assign  image_0_106[39:32]   = Image[145];
    assign  image_0_106[31:24]   = Image[146];
    assign  image_0_106[23:16]   = Image[176];
    assign  image_0_106[15:8]    = Image[177];
    assign  image_0_106[7:0]     = Image[178];

    assign  image_0_107[71:64]   = Image[113];
    assign  image_0_107[63:56]   = Image[114];
    assign  image_0_107[55:48]   = Image[115];
    assign  image_0_107[47:40]   = Image[145];
    assign  image_0_107[39:32]   = Image[146];
    assign  image_0_107[31:24]   = Image[147];
    assign  image_0_107[23:16]   = Image[177];
    assign  image_0_107[15:8]    = Image[178];
    assign  image_0_107[7:0]     = Image[179];

    assign  image_0_108[71:64]   = Image[114];
    assign  image_0_108[63:56]   = Image[115];
    assign  image_0_108[55:48]   = Image[116];
    assign  image_0_108[47:40]   = Image[146];
    assign  image_0_108[39:32]   = Image[147];
    assign  image_0_108[31:24]   = Image[148];
    assign  image_0_108[23:16]   = Image[178];
    assign  image_0_108[15:8]    = Image[179];
    assign  image_0_108[7:0]     = Image[180];

    assign  image_0_109[71:64]   = Image[115];
    assign  image_0_109[63:56]   = Image[116];
    assign  image_0_109[55:48]   = Image[117];
    assign  image_0_109[47:40]   = Image[147];
    assign  image_0_109[39:32]   = Image[148];
    assign  image_0_109[31:24]   = Image[149];
    assign  image_0_109[23:16]   = Image[179];
    assign  image_0_109[15:8]    = Image[180];
    assign  image_0_109[7:0]     = Image[181];

    assign  image_0_110[71:64]   = Image[116];
    assign  image_0_110[63:56]   = Image[117];
    assign  image_0_110[55:48]   = Image[118];
    assign  image_0_110[47:40]   = Image[148];
    assign  image_0_110[39:32]   = Image[149];
    assign  image_0_110[31:24]   = Image[150];
    assign  image_0_110[23:16]   = Image[180];
    assign  image_0_110[15:8]    = Image[181];
    assign  image_0_110[7:0]     = Image[182];

    assign  image_0_111[71:64]   = Image[117];
    assign  image_0_111[63:56]   = Image[118];
    assign  image_0_111[55:48]   = Image[119];
    assign  image_0_111[47:40]   = Image[149];
    assign  image_0_111[39:32]   = Image[150];
    assign  image_0_111[31:24]   = Image[151];
    assign  image_0_111[23:16]   = Image[181];
    assign  image_0_111[15:8]    = Image[182];
    assign  image_0_111[7:0]     = Image[183];

    assign  image_0_112[71:64]   = Image[118];
    assign  image_0_112[63:56]   = Image[119];
    assign  image_0_112[55:48]   = Image[120];
    assign  image_0_112[47:40]   = Image[150];
    assign  image_0_112[39:32]   = Image[151];
    assign  image_0_112[31:24]   = Image[152];
    assign  image_0_112[23:16]   = Image[182];
    assign  image_0_112[15:8]    = Image[183];
    assign  image_0_112[7:0]     = Image[184];

    assign  image_0_113[71:64]   = Image[119];
    assign  image_0_113[63:56]   = Image[120];
    assign  image_0_113[55:48]   = Image[121];
    assign  image_0_113[47:40]   = Image[151];
    assign  image_0_113[39:32]   = Image[152];
    assign  image_0_113[31:24]   = Image[153];
    assign  image_0_113[23:16]   = Image[183];
    assign  image_0_113[15:8]    = Image[184];
    assign  image_0_113[7:0]     = Image[185];

    assign  image_0_114[71:64]   = Image[120];
    assign  image_0_114[63:56]   = Image[121];
    assign  image_0_114[55:48]   = Image[122];
    assign  image_0_114[47:40]   = Image[152];
    assign  image_0_114[39:32]   = Image[153];
    assign  image_0_114[31:24]   = Image[154];
    assign  image_0_114[23:16]   = Image[184];
    assign  image_0_114[15:8]    = Image[185];
    assign  image_0_114[7:0]     = Image[186];

    assign  image_0_115[71:64]   = Image[121];
    assign  image_0_115[63:56]   = Image[122];
    assign  image_0_115[55:48]   = Image[123];
    assign  image_0_115[47:40]   = Image[153];
    assign  image_0_115[39:32]   = Image[154];
    assign  image_0_115[31:24]   = Image[155];
    assign  image_0_115[23:16]   = Image[185];
    assign  image_0_115[15:8]    = Image[186];
    assign  image_0_115[7:0]     = Image[187];

    assign  image_0_116[71:64]   = Image[122];
    assign  image_0_116[63:56]   = Image[123];
    assign  image_0_116[55:48]   = Image[124];
    assign  image_0_116[47:40]   = Image[154];
    assign  image_0_116[39:32]   = Image[155];
    assign  image_0_116[31:24]   = Image[156];
    assign  image_0_116[23:16]   = Image[186];
    assign  image_0_116[15:8]    = Image[187];
    assign  image_0_116[7:0]     = Image[188];

    assign  image_0_117[71:64]   = Image[123];
    assign  image_0_117[63:56]   = Image[124];
    assign  image_0_117[55:48]   = Image[125];
    assign  image_0_117[47:40]   = Image[155];
    assign  image_0_117[39:32]   = Image[156];
    assign  image_0_117[31:24]   = Image[157];
    assign  image_0_117[23:16]   = Image[187];
    assign  image_0_117[15:8]    = Image[188];
    assign  image_0_117[7:0]     = Image[189];

    assign  image_0_118[71:64]   = Image[124];
    assign  image_0_118[63:56]   = Image[125];
    assign  image_0_118[55:48]   = Image[126];
    assign  image_0_118[47:40]   = Image[156];
    assign  image_0_118[39:32]   = Image[157];
    assign  image_0_118[31:24]   = Image[158];
    assign  image_0_118[23:16]   = Image[188];
    assign  image_0_118[15:8]    = Image[189];
    assign  image_0_118[7:0]     = Image[190];

    assign  image_0_119[71:64]   = Image[125];
    assign  image_0_119[63:56]   = Image[126];
    assign  image_0_119[55:48]   = Image[127];
    assign  image_0_119[47:40]   = Image[157];
    assign  image_0_119[39:32]   = Image[158];
    assign  image_0_119[31:24]   = Image[159];
    assign  image_0_119[23:16]   = Image[189];
    assign  image_0_119[15:8]    = Image[190];
    assign  image_0_119[7:0]     = Image[191];

    assign  image_0_120[71:64]   = Image[128];
    assign  image_0_120[63:56]   = Image[129];
    assign  image_0_120[55:48]   = Image[130];
    assign  image_0_120[47:40]   = Image[160];
    assign  image_0_120[39:32]   = Image[161];
    assign  image_0_120[31:24]   = Image[162];
    assign  image_0_120[23:16]   = Image[192];
    assign  image_0_120[15:8]    = Image[193];
    assign  image_0_120[7:0]     = Image[194];

    assign  image_0_121[71:64]   = Image[129];
    assign  image_0_121[63:56]   = Image[130];
    assign  image_0_121[55:48]   = Image[131];
    assign  image_0_121[47:40]   = Image[161];
    assign  image_0_121[39:32]   = Image[162];
    assign  image_0_121[31:24]   = Image[163];
    assign  image_0_121[23:16]   = Image[193];
    assign  image_0_121[15:8]    = Image[194];
    assign  image_0_121[7:0]     = Image[195];

    assign  image_0_122[71:64]   = Image[130];
    assign  image_0_122[63:56]   = Image[131];
    assign  image_0_122[55:48]   = Image[132];
    assign  image_0_122[47:40]   = Image[162];
    assign  image_0_122[39:32]   = Image[163];
    assign  image_0_122[31:24]   = Image[164];
    assign  image_0_122[23:16]   = Image[194];
    assign  image_0_122[15:8]    = Image[195];
    assign  image_0_122[7:0]     = Image[196];

    assign  image_0_123[71:64]   = Image[131];
    assign  image_0_123[63:56]   = Image[132];
    assign  image_0_123[55:48]   = Image[133];
    assign  image_0_123[47:40]   = Image[163];
    assign  image_0_123[39:32]   = Image[164];
    assign  image_0_123[31:24]   = Image[165];
    assign  image_0_123[23:16]   = Image[195];
    assign  image_0_123[15:8]    = Image[196];
    assign  image_0_123[7:0]     = Image[197];

    assign  image_0_124[71:64]   = Image[132];
    assign  image_0_124[63:56]   = Image[133];
    assign  image_0_124[55:48]   = Image[134];
    assign  image_0_124[47:40]   = Image[164];
    assign  image_0_124[39:32]   = Image[165];
    assign  image_0_124[31:24]   = Image[166];
    assign  image_0_124[23:16]   = Image[196];
    assign  image_0_124[15:8]    = Image[197];
    assign  image_0_124[7:0]     = Image[198];

    assign  image_0_125[71:64]   = Image[133];
    assign  image_0_125[63:56]   = Image[134];
    assign  image_0_125[55:48]   = Image[135];
    assign  image_0_125[47:40]   = Image[165];
    assign  image_0_125[39:32]   = Image[166];
    assign  image_0_125[31:24]   = Image[167];
    assign  image_0_125[23:16]   = Image[197];
    assign  image_0_125[15:8]    = Image[198];
    assign  image_0_125[7:0]     = Image[199];

    assign  image_0_126[71:64]   = Image[134];
    assign  image_0_126[63:56]   = Image[135];
    assign  image_0_126[55:48]   = Image[136];
    assign  image_0_126[47:40]   = Image[166];
    assign  image_0_126[39:32]   = Image[167];
    assign  image_0_126[31:24]   = Image[168];
    assign  image_0_126[23:16]   = Image[198];
    assign  image_0_126[15:8]    = Image[199];
    assign  image_0_126[7:0]     = Image[200];

    assign  image_0_127[71:64]   = Image[135];
    assign  image_0_127[63:56]   = Image[136];
    assign  image_0_127[55:48]   = Image[137];
    assign  image_0_127[47:40]   = Image[167];
    assign  image_0_127[39:32]   = Image[168];
    assign  image_0_127[31:24]   = Image[169];
    assign  image_0_127[23:16]   = Image[199];
    assign  image_0_127[15:8]    = Image[200];
    assign  image_0_127[7:0]     = Image[201];

    assign  image_0_128[71:64]   = Image[136];
    assign  image_0_128[63:56]   = Image[137];
    assign  image_0_128[55:48]   = Image[138];
    assign  image_0_128[47:40]   = Image[168];
    assign  image_0_128[39:32]   = Image[169];
    assign  image_0_128[31:24]   = Image[170];
    assign  image_0_128[23:16]   = Image[200];
    assign  image_0_128[15:8]    = Image[201];
    assign  image_0_128[7:0]     = Image[202];

    assign  image_0_129[71:64]   = Image[137];
    assign  image_0_129[63:56]   = Image[138];
    assign  image_0_129[55:48]   = Image[139];
    assign  image_0_129[47:40]   = Image[169];
    assign  image_0_129[39:32]   = Image[170];
    assign  image_0_129[31:24]   = Image[171];
    assign  image_0_129[23:16]   = Image[201];
    assign  image_0_129[15:8]    = Image[202];
    assign  image_0_129[7:0]     = Image[203];

    assign  image_0_130[71:64]   = Image[138];
    assign  image_0_130[63:56]   = Image[139];
    assign  image_0_130[55:48]   = Image[140];
    assign  image_0_130[47:40]   = Image[170];
    assign  image_0_130[39:32]   = Image[171];
    assign  image_0_130[31:24]   = Image[172];
    assign  image_0_130[23:16]   = Image[202];
    assign  image_0_130[15:8]    = Image[203];
    assign  image_0_130[7:0]     = Image[204];

    assign  image_0_131[71:64]   = Image[139];
    assign  image_0_131[63:56]   = Image[140];
    assign  image_0_131[55:48]   = Image[141];
    assign  image_0_131[47:40]   = Image[171];
    assign  image_0_131[39:32]   = Image[172];
    assign  image_0_131[31:24]   = Image[173];
    assign  image_0_131[23:16]   = Image[203];
    assign  image_0_131[15:8]    = Image[204];
    assign  image_0_131[7:0]     = Image[205];

    assign  image_0_132[71:64]   = Image[140];
    assign  image_0_132[63:56]   = Image[141];
    assign  image_0_132[55:48]   = Image[142];
    assign  image_0_132[47:40]   = Image[172];
    assign  image_0_132[39:32]   = Image[173];
    assign  image_0_132[31:24]   = Image[174];
    assign  image_0_132[23:16]   = Image[204];
    assign  image_0_132[15:8]    = Image[205];
    assign  image_0_132[7:0]     = Image[206];

    assign  image_0_133[71:64]   = Image[141];
    assign  image_0_133[63:56]   = Image[142];
    assign  image_0_133[55:48]   = Image[143];
    assign  image_0_133[47:40]   = Image[173];
    assign  image_0_133[39:32]   = Image[174];
    assign  image_0_133[31:24]   = Image[175];
    assign  image_0_133[23:16]   = Image[205];
    assign  image_0_133[15:8]    = Image[206];
    assign  image_0_133[7:0]     = Image[207];

    assign  image_0_134[71:64]   = Image[142];
    assign  image_0_134[63:56]   = Image[143];
    assign  image_0_134[55:48]   = Image[144];
    assign  image_0_134[47:40]   = Image[174];
    assign  image_0_134[39:32]   = Image[175];
    assign  image_0_134[31:24]   = Image[176];
    assign  image_0_134[23:16]   = Image[206];
    assign  image_0_134[15:8]    = Image[207];
    assign  image_0_134[7:0]     = Image[208];

    assign  image_0_135[71:64]   = Image[143];
    assign  image_0_135[63:56]   = Image[144];
    assign  image_0_135[55:48]   = Image[145];
    assign  image_0_135[47:40]   = Image[175];
    assign  image_0_135[39:32]   = Image[176];
    assign  image_0_135[31:24]   = Image[177];
    assign  image_0_135[23:16]   = Image[207];
    assign  image_0_135[15:8]    = Image[208];
    assign  image_0_135[7:0]     = Image[209];

    assign  image_0_136[71:64]   = Image[144];
    assign  image_0_136[63:56]   = Image[145];
    assign  image_0_136[55:48]   = Image[146];
    assign  image_0_136[47:40]   = Image[176];
    assign  image_0_136[39:32]   = Image[177];
    assign  image_0_136[31:24]   = Image[178];
    assign  image_0_136[23:16]   = Image[208];
    assign  image_0_136[15:8]    = Image[209];
    assign  image_0_136[7:0]     = Image[210];

    assign  image_0_137[71:64]   = Image[145];
    assign  image_0_137[63:56]   = Image[146];
    assign  image_0_137[55:48]   = Image[147];
    assign  image_0_137[47:40]   = Image[177];
    assign  image_0_137[39:32]   = Image[178];
    assign  image_0_137[31:24]   = Image[179];
    assign  image_0_137[23:16]   = Image[209];
    assign  image_0_137[15:8]    = Image[210];
    assign  image_0_137[7:0]     = Image[211];

    assign  image_0_138[71:64]   = Image[146];
    assign  image_0_138[63:56]   = Image[147];
    assign  image_0_138[55:48]   = Image[148];
    assign  image_0_138[47:40]   = Image[178];
    assign  image_0_138[39:32]   = Image[179];
    assign  image_0_138[31:24]   = Image[180];
    assign  image_0_138[23:16]   = Image[210];
    assign  image_0_138[15:8]    = Image[211];
    assign  image_0_138[7:0]     = Image[212];

    assign  image_0_139[71:64]   = Image[147];
    assign  image_0_139[63:56]   = Image[148];
    assign  image_0_139[55:48]   = Image[149];
    assign  image_0_139[47:40]   = Image[179];
    assign  image_0_139[39:32]   = Image[180];
    assign  image_0_139[31:24]   = Image[181];
    assign  image_0_139[23:16]   = Image[211];
    assign  image_0_139[15:8]    = Image[212];
    assign  image_0_139[7:0]     = Image[213];

    assign  image_0_140[71:64]   = Image[148];
    assign  image_0_140[63:56]   = Image[149];
    assign  image_0_140[55:48]   = Image[150];
    assign  image_0_140[47:40]   = Image[180];
    assign  image_0_140[39:32]   = Image[181];
    assign  image_0_140[31:24]   = Image[182];
    assign  image_0_140[23:16]   = Image[212];
    assign  image_0_140[15:8]    = Image[213];
    assign  image_0_140[7:0]     = Image[214];

    assign  image_0_141[71:64]   = Image[149];
    assign  image_0_141[63:56]   = Image[150];
    assign  image_0_141[55:48]   = Image[151];
    assign  image_0_141[47:40]   = Image[181];
    assign  image_0_141[39:32]   = Image[182];
    assign  image_0_141[31:24]   = Image[183];
    assign  image_0_141[23:16]   = Image[213];
    assign  image_0_141[15:8]    = Image[214];
    assign  image_0_141[7:0]     = Image[215];

    assign  image_0_142[71:64]   = Image[150];
    assign  image_0_142[63:56]   = Image[151];
    assign  image_0_142[55:48]   = Image[152];
    assign  image_0_142[47:40]   = Image[182];
    assign  image_0_142[39:32]   = Image[183];
    assign  image_0_142[31:24]   = Image[184];
    assign  image_0_142[23:16]   = Image[214];
    assign  image_0_142[15:8]    = Image[215];
    assign  image_0_142[7:0]     = Image[216];

    assign  image_0_143[71:64]   = Image[151];
    assign  image_0_143[63:56]   = Image[152];
    assign  image_0_143[55:48]   = Image[153];
    assign  image_0_143[47:40]   = Image[183];
    assign  image_0_143[39:32]   = Image[184];
    assign  image_0_143[31:24]   = Image[185];
    assign  image_0_143[23:16]   = Image[215];
    assign  image_0_143[15:8]    = Image[216];
    assign  image_0_143[7:0]     = Image[217];

    assign  image_0_144[71:64]   = Image[152];
    assign  image_0_144[63:56]   = Image[153];
    assign  image_0_144[55:48]   = Image[154];
    assign  image_0_144[47:40]   = Image[184];
    assign  image_0_144[39:32]   = Image[185];
    assign  image_0_144[31:24]   = Image[186];
    assign  image_0_144[23:16]   = Image[216];
    assign  image_0_144[15:8]    = Image[217];
    assign  image_0_144[7:0]     = Image[218];

    assign  image_0_145[71:64]   = Image[153];
    assign  image_0_145[63:56]   = Image[154];
    assign  image_0_145[55:48]   = Image[155];
    assign  image_0_145[47:40]   = Image[185];
    assign  image_0_145[39:32]   = Image[186];
    assign  image_0_145[31:24]   = Image[187];
    assign  image_0_145[23:16]   = Image[217];
    assign  image_0_145[15:8]    = Image[218];
    assign  image_0_145[7:0]     = Image[219];

    assign  image_0_146[71:64]   = Image[154];
    assign  image_0_146[63:56]   = Image[155];
    assign  image_0_146[55:48]   = Image[156];
    assign  image_0_146[47:40]   = Image[186];
    assign  image_0_146[39:32]   = Image[187];
    assign  image_0_146[31:24]   = Image[188];
    assign  image_0_146[23:16]   = Image[218];
    assign  image_0_146[15:8]    = Image[219];
    assign  image_0_146[7:0]     = Image[220];

    assign  image_0_147[71:64]   = Image[155];
    assign  image_0_147[63:56]   = Image[156];
    assign  image_0_147[55:48]   = Image[157];
    assign  image_0_147[47:40]   = Image[187];
    assign  image_0_147[39:32]   = Image[188];
    assign  image_0_147[31:24]   = Image[189];
    assign  image_0_147[23:16]   = Image[219];
    assign  image_0_147[15:8]    = Image[220];
    assign  image_0_147[7:0]     = Image[221];

    assign  image_0_148[71:64]   = Image[156];
    assign  image_0_148[63:56]   = Image[157];
    assign  image_0_148[55:48]   = Image[158];
    assign  image_0_148[47:40]   = Image[188];
    assign  image_0_148[39:32]   = Image[189];
    assign  image_0_148[31:24]   = Image[190];
    assign  image_0_148[23:16]   = Image[220];
    assign  image_0_148[15:8]    = Image[221];
    assign  image_0_148[7:0]     = Image[222];

    assign  image_0_149[71:64]   = Image[157];
    assign  image_0_149[63:56]   = Image[158];
    assign  image_0_149[55:48]   = Image[159];
    assign  image_0_149[47:40]   = Image[189];
    assign  image_0_149[39:32]   = Image[190];
    assign  image_0_149[31:24]   = Image[191];
    assign  image_0_149[23:16]   = Image[221];
    assign  image_0_149[15:8]    = Image[222];
    assign  image_0_149[7:0]     = Image[223];

    assign  image_0_150[71:64]   = Image[160];
    assign  image_0_150[63:56]   = Image[161];
    assign  image_0_150[55:48]   = Image[162];
    assign  image_0_150[47:40]   = Image[192];
    assign  image_0_150[39:32]   = Image[193];
    assign  image_0_150[31:24]   = Image[194];
    assign  image_0_150[23:16]   = Image[224];
    assign  image_0_150[15:8]    = Image[225];
    assign  image_0_150[7:0]     = Image[226];

    assign  image_0_151[71:64]   = Image[161];
    assign  image_0_151[63:56]   = Image[162];
    assign  image_0_151[55:48]   = Image[163];
    assign  image_0_151[47:40]   = Image[193];
    assign  image_0_151[39:32]   = Image[194];
    assign  image_0_151[31:24]   = Image[195];
    assign  image_0_151[23:16]   = Image[225];
    assign  image_0_151[15:8]    = Image[226];
    assign  image_0_151[7:0]     = Image[227];

    assign  image_0_152[71:64]   = Image[162];
    assign  image_0_152[63:56]   = Image[163];
    assign  image_0_152[55:48]   = Image[164];
    assign  image_0_152[47:40]   = Image[194];
    assign  image_0_152[39:32]   = Image[195];
    assign  image_0_152[31:24]   = Image[196];
    assign  image_0_152[23:16]   = Image[226];
    assign  image_0_152[15:8]    = Image[227];
    assign  image_0_152[7:0]     = Image[228];

    assign  image_0_153[71:64]   = Image[163];
    assign  image_0_153[63:56]   = Image[164];
    assign  image_0_153[55:48]   = Image[165];
    assign  image_0_153[47:40]   = Image[195];
    assign  image_0_153[39:32]   = Image[196];
    assign  image_0_153[31:24]   = Image[197];
    assign  image_0_153[23:16]   = Image[227];
    assign  image_0_153[15:8]    = Image[228];
    assign  image_0_153[7:0]     = Image[229];

    assign  image_0_154[71:64]   = Image[164];
    assign  image_0_154[63:56]   = Image[165];
    assign  image_0_154[55:48]   = Image[166];
    assign  image_0_154[47:40]   = Image[196];
    assign  image_0_154[39:32]   = Image[197];
    assign  image_0_154[31:24]   = Image[198];
    assign  image_0_154[23:16]   = Image[228];
    assign  image_0_154[15:8]    = Image[229];
    assign  image_0_154[7:0]     = Image[230];

    assign  image_0_155[71:64]   = Image[165];
    assign  image_0_155[63:56]   = Image[166];
    assign  image_0_155[55:48]   = Image[167];
    assign  image_0_155[47:40]   = Image[197];
    assign  image_0_155[39:32]   = Image[198];
    assign  image_0_155[31:24]   = Image[199];
    assign  image_0_155[23:16]   = Image[229];
    assign  image_0_155[15:8]    = Image[230];
    assign  image_0_155[7:0]     = Image[231];

    assign  image_0_156[71:64]   = Image[166];
    assign  image_0_156[63:56]   = Image[167];
    assign  image_0_156[55:48]   = Image[168];
    assign  image_0_156[47:40]   = Image[198];
    assign  image_0_156[39:32]   = Image[199];
    assign  image_0_156[31:24]   = Image[200];
    assign  image_0_156[23:16]   = Image[230];
    assign  image_0_156[15:8]    = Image[231];
    assign  image_0_156[7:0]     = Image[232];

    assign  image_0_157[71:64]   = Image[167];
    assign  image_0_157[63:56]   = Image[168];
    assign  image_0_157[55:48]   = Image[169];
    assign  image_0_157[47:40]   = Image[199];
    assign  image_0_157[39:32]   = Image[200];
    assign  image_0_157[31:24]   = Image[201];
    assign  image_0_157[23:16]   = Image[231];
    assign  image_0_157[15:8]    = Image[232];
    assign  image_0_157[7:0]     = Image[233];

    assign  image_0_158[71:64]   = Image[168];
    assign  image_0_158[63:56]   = Image[169];
    assign  image_0_158[55:48]   = Image[170];
    assign  image_0_158[47:40]   = Image[200];
    assign  image_0_158[39:32]   = Image[201];
    assign  image_0_158[31:24]   = Image[202];
    assign  image_0_158[23:16]   = Image[232];
    assign  image_0_158[15:8]    = Image[233];
    assign  image_0_158[7:0]     = Image[234];

    assign  image_0_159[71:64]   = Image[169];
    assign  image_0_159[63:56]   = Image[170];
    assign  image_0_159[55:48]   = Image[171];
    assign  image_0_159[47:40]   = Image[201];
    assign  image_0_159[39:32]   = Image[202];
    assign  image_0_159[31:24]   = Image[203];
    assign  image_0_159[23:16]   = Image[233];
    assign  image_0_159[15:8]    = Image[234];
    assign  image_0_159[7:0]     = Image[235];

    assign  image_0_160[71:64]   = Image[170];
    assign  image_0_160[63:56]   = Image[171];
    assign  image_0_160[55:48]   = Image[172];
    assign  image_0_160[47:40]   = Image[202];
    assign  image_0_160[39:32]   = Image[203];
    assign  image_0_160[31:24]   = Image[204];
    assign  image_0_160[23:16]   = Image[234];
    assign  image_0_160[15:8]    = Image[235];
    assign  image_0_160[7:0]     = Image[236];

    assign  image_0_161[71:64]   = Image[171];
    assign  image_0_161[63:56]   = Image[172];
    assign  image_0_161[55:48]   = Image[173];
    assign  image_0_161[47:40]   = Image[203];
    assign  image_0_161[39:32]   = Image[204];
    assign  image_0_161[31:24]   = Image[205];
    assign  image_0_161[23:16]   = Image[235];
    assign  image_0_161[15:8]    = Image[236];
    assign  image_0_161[7:0]     = Image[237];

    assign  image_0_162[71:64]   = Image[172];
    assign  image_0_162[63:56]   = Image[173];
    assign  image_0_162[55:48]   = Image[174];
    assign  image_0_162[47:40]   = Image[204];
    assign  image_0_162[39:32]   = Image[205];
    assign  image_0_162[31:24]   = Image[206];
    assign  image_0_162[23:16]   = Image[236];
    assign  image_0_162[15:8]    = Image[237];
    assign  image_0_162[7:0]     = Image[238];

    assign  image_0_163[71:64]   = Image[173];
    assign  image_0_163[63:56]   = Image[174];
    assign  image_0_163[55:48]   = Image[175];
    assign  image_0_163[47:40]   = Image[205];
    assign  image_0_163[39:32]   = Image[206];
    assign  image_0_163[31:24]   = Image[207];
    assign  image_0_163[23:16]   = Image[237];
    assign  image_0_163[15:8]    = Image[238];
    assign  image_0_163[7:0]     = Image[239];

    assign  image_0_164[71:64]   = Image[174];
    assign  image_0_164[63:56]   = Image[175];
    assign  image_0_164[55:48]   = Image[176];
    assign  image_0_164[47:40]   = Image[206];
    assign  image_0_164[39:32]   = Image[207];
    assign  image_0_164[31:24]   = Image[208];
    assign  image_0_164[23:16]   = Image[238];
    assign  image_0_164[15:8]    = Image[239];
    assign  image_0_164[7:0]     = Image[240];

    assign  image_0_165[71:64]   = Image[175];
    assign  image_0_165[63:56]   = Image[176];
    assign  image_0_165[55:48]   = Image[177];
    assign  image_0_165[47:40]   = Image[207];
    assign  image_0_165[39:32]   = Image[208];
    assign  image_0_165[31:24]   = Image[209];
    assign  image_0_165[23:16]   = Image[239];
    assign  image_0_165[15:8]    = Image[240];
    assign  image_0_165[7:0]     = Image[241];

    assign  image_0_166[71:64]   = Image[176];
    assign  image_0_166[63:56]   = Image[177];
    assign  image_0_166[55:48]   = Image[178];
    assign  image_0_166[47:40]   = Image[208];
    assign  image_0_166[39:32]   = Image[209];
    assign  image_0_166[31:24]   = Image[210];
    assign  image_0_166[23:16]   = Image[240];
    assign  image_0_166[15:8]    = Image[241];
    assign  image_0_166[7:0]     = Image[242];

    assign  image_0_167[71:64]   = Image[177];
    assign  image_0_167[63:56]   = Image[178];
    assign  image_0_167[55:48]   = Image[179];
    assign  image_0_167[47:40]   = Image[209];
    assign  image_0_167[39:32]   = Image[210];
    assign  image_0_167[31:24]   = Image[211];
    assign  image_0_167[23:16]   = Image[241];
    assign  image_0_167[15:8]    = Image[242];
    assign  image_0_167[7:0]     = Image[243];

    assign  image_0_168[71:64]   = Image[178];
    assign  image_0_168[63:56]   = Image[179];
    assign  image_0_168[55:48]   = Image[180];
    assign  image_0_168[47:40]   = Image[210];
    assign  image_0_168[39:32]   = Image[211];
    assign  image_0_168[31:24]   = Image[212];
    assign  image_0_168[23:16]   = Image[242];
    assign  image_0_168[15:8]    = Image[243];
    assign  image_0_168[7:0]     = Image[244];

    assign  image_0_169[71:64]   = Image[179];
    assign  image_0_169[63:56]   = Image[180];
    assign  image_0_169[55:48]   = Image[181];
    assign  image_0_169[47:40]   = Image[211];
    assign  image_0_169[39:32]   = Image[212];
    assign  image_0_169[31:24]   = Image[213];
    assign  image_0_169[23:16]   = Image[243];
    assign  image_0_169[15:8]    = Image[244];
    assign  image_0_169[7:0]     = Image[245];

    assign  image_0_170[71:64]   = Image[180];
    assign  image_0_170[63:56]   = Image[181];
    assign  image_0_170[55:48]   = Image[182];
    assign  image_0_170[47:40]   = Image[212];
    assign  image_0_170[39:32]   = Image[213];
    assign  image_0_170[31:24]   = Image[214];
    assign  image_0_170[23:16]   = Image[244];
    assign  image_0_170[15:8]    = Image[245];
    assign  image_0_170[7:0]     = Image[246];

    assign  image_0_171[71:64]   = Image[181];
    assign  image_0_171[63:56]   = Image[182];
    assign  image_0_171[55:48]   = Image[183];
    assign  image_0_171[47:40]   = Image[213];
    assign  image_0_171[39:32]   = Image[214];
    assign  image_0_171[31:24]   = Image[215];
    assign  image_0_171[23:16]   = Image[245];
    assign  image_0_171[15:8]    = Image[246];
    assign  image_0_171[7:0]     = Image[247];

    assign  image_0_172[71:64]   = Image[182];
    assign  image_0_172[63:56]   = Image[183];
    assign  image_0_172[55:48]   = Image[184];
    assign  image_0_172[47:40]   = Image[214];
    assign  image_0_172[39:32]   = Image[215];
    assign  image_0_172[31:24]   = Image[216];
    assign  image_0_172[23:16]   = Image[246];
    assign  image_0_172[15:8]    = Image[247];
    assign  image_0_172[7:0]     = Image[248];

    assign  image_0_173[71:64]   = Image[183];
    assign  image_0_173[63:56]   = Image[184];
    assign  image_0_173[55:48]   = Image[185];
    assign  image_0_173[47:40]   = Image[215];
    assign  image_0_173[39:32]   = Image[216];
    assign  image_0_173[31:24]   = Image[217];
    assign  image_0_173[23:16]   = Image[247];
    assign  image_0_173[15:8]    = Image[248];
    assign  image_0_173[7:0]     = Image[249];

    assign  image_0_174[71:64]   = Image[184];
    assign  image_0_174[63:56]   = Image[185];
    assign  image_0_174[55:48]   = Image[186];
    assign  image_0_174[47:40]   = Image[216];
    assign  image_0_174[39:32]   = Image[217];
    assign  image_0_174[31:24]   = Image[218];
    assign  image_0_174[23:16]   = Image[248];
    assign  image_0_174[15:8]    = Image[249];
    assign  image_0_174[7:0]     = Image[250];

    assign  image_0_175[71:64]   = Image[185];
    assign  image_0_175[63:56]   = Image[186];
    assign  image_0_175[55:48]   = Image[187];
    assign  image_0_175[47:40]   = Image[217];
    assign  image_0_175[39:32]   = Image[218];
    assign  image_0_175[31:24]   = Image[219];
    assign  image_0_175[23:16]   = Image[249];
    assign  image_0_175[15:8]    = Image[250];
    assign  image_0_175[7:0]     = Image[251];

    assign  image_0_176[71:64]   = Image[186];
    assign  image_0_176[63:56]   = Image[187];
    assign  image_0_176[55:48]   = Image[188];
    assign  image_0_176[47:40]   = Image[218];
    assign  image_0_176[39:32]   = Image[219];
    assign  image_0_176[31:24]   = Image[220];
    assign  image_0_176[23:16]   = Image[250];
    assign  image_0_176[15:8]    = Image[251];
    assign  image_0_176[7:0]     = Image[252];

    assign  image_0_177[71:64]   = Image[187];
    assign  image_0_177[63:56]   = Image[188];
    assign  image_0_177[55:48]   = Image[189];
    assign  image_0_177[47:40]   = Image[219];
    assign  image_0_177[39:32]   = Image[220];
    assign  image_0_177[31:24]   = Image[221];
    assign  image_0_177[23:16]   = Image[251];
    assign  image_0_177[15:8]    = Image[252];
    assign  image_0_177[7:0]     = Image[253];

    assign  image_0_178[71:64]   = Image[188];
    assign  image_0_178[63:56]   = Image[189];
    assign  image_0_178[55:48]   = Image[190];
    assign  image_0_178[47:40]   = Image[220];
    assign  image_0_178[39:32]   = Image[221];
    assign  image_0_178[31:24]   = Image[222];
    assign  image_0_178[23:16]   = Image[252];
    assign  image_0_178[15:8]    = Image[253];
    assign  image_0_178[7:0]     = Image[254];

    assign  image_0_179[71:64]   = Image[189];
    assign  image_0_179[63:56]   = Image[190];
    assign  image_0_179[55:48]   = Image[191];
    assign  image_0_179[47:40]   = Image[221];
    assign  image_0_179[39:32]   = Image[222];
    assign  image_0_179[31:24]   = Image[223];
    assign  image_0_179[23:16]   = Image[253];
    assign  image_0_179[15:8]    = Image[254];
    assign  image_0_179[7:0]     = Image[255];

    assign  image_0_180[71:64]   = Image[192];
    assign  image_0_180[63:56]   = Image[193];
    assign  image_0_180[55:48]   = Image[194];
    assign  image_0_180[47:40]   = Image[224];
    assign  image_0_180[39:32]   = Image[225];
    assign  image_0_180[31:24]   = Image[226];
    assign  image_0_180[23:16]   = Image[256];
    assign  image_0_180[15:8]    = Image[257];
    assign  image_0_180[7:0]     = Image[258];

    assign  image_0_181[71:64]   = Image[193];
    assign  image_0_181[63:56]   = Image[194];
    assign  image_0_181[55:48]   = Image[195];
    assign  image_0_181[47:40]   = Image[225];
    assign  image_0_181[39:32]   = Image[226];
    assign  image_0_181[31:24]   = Image[227];
    assign  image_0_181[23:16]   = Image[257];
    assign  image_0_181[15:8]    = Image[258];
    assign  image_0_181[7:0]     = Image[259];

    assign  image_0_182[71:64]   = Image[194];
    assign  image_0_182[63:56]   = Image[195];
    assign  image_0_182[55:48]   = Image[196];
    assign  image_0_182[47:40]   = Image[226];
    assign  image_0_182[39:32]   = Image[227];
    assign  image_0_182[31:24]   = Image[228];
    assign  image_0_182[23:16]   = Image[258];
    assign  image_0_182[15:8]    = Image[259];
    assign  image_0_182[7:0]     = Image[260];

    assign  image_0_183[71:64]   = Image[195];
    assign  image_0_183[63:56]   = Image[196];
    assign  image_0_183[55:48]   = Image[197];
    assign  image_0_183[47:40]   = Image[227];
    assign  image_0_183[39:32]   = Image[228];
    assign  image_0_183[31:24]   = Image[229];
    assign  image_0_183[23:16]   = Image[259];
    assign  image_0_183[15:8]    = Image[260];
    assign  image_0_183[7:0]     = Image[261];

    assign  image_0_184[71:64]   = Image[196];
    assign  image_0_184[63:56]   = Image[197];
    assign  image_0_184[55:48]   = Image[198];
    assign  image_0_184[47:40]   = Image[228];
    assign  image_0_184[39:32]   = Image[229];
    assign  image_0_184[31:24]   = Image[230];
    assign  image_0_184[23:16]   = Image[260];
    assign  image_0_184[15:8]    = Image[261];
    assign  image_0_184[7:0]     = Image[262];

    assign  image_0_185[71:64]   = Image[197];
    assign  image_0_185[63:56]   = Image[198];
    assign  image_0_185[55:48]   = Image[199];
    assign  image_0_185[47:40]   = Image[229];
    assign  image_0_185[39:32]   = Image[230];
    assign  image_0_185[31:24]   = Image[231];
    assign  image_0_185[23:16]   = Image[261];
    assign  image_0_185[15:8]    = Image[262];
    assign  image_0_185[7:0]     = Image[263];

    assign  image_0_186[71:64]   = Image[198];
    assign  image_0_186[63:56]   = Image[199];
    assign  image_0_186[55:48]   = Image[200];
    assign  image_0_186[47:40]   = Image[230];
    assign  image_0_186[39:32]   = Image[231];
    assign  image_0_186[31:24]   = Image[232];
    assign  image_0_186[23:16]   = Image[262];
    assign  image_0_186[15:8]    = Image[263];
    assign  image_0_186[7:0]     = Image[264];

    assign  image_0_187[71:64]   = Image[199];
    assign  image_0_187[63:56]   = Image[200];
    assign  image_0_187[55:48]   = Image[201];
    assign  image_0_187[47:40]   = Image[231];
    assign  image_0_187[39:32]   = Image[232];
    assign  image_0_187[31:24]   = Image[233];
    assign  image_0_187[23:16]   = Image[263];
    assign  image_0_187[15:8]    = Image[264];
    assign  image_0_187[7:0]     = Image[265];

    assign  image_0_188[71:64]   = Image[200];
    assign  image_0_188[63:56]   = Image[201];
    assign  image_0_188[55:48]   = Image[202];
    assign  image_0_188[47:40]   = Image[232];
    assign  image_0_188[39:32]   = Image[233];
    assign  image_0_188[31:24]   = Image[234];
    assign  image_0_188[23:16]   = Image[264];
    assign  image_0_188[15:8]    = Image[265];
    assign  image_0_188[7:0]     = Image[266];

    assign  image_0_189[71:64]   = Image[201];
    assign  image_0_189[63:56]   = Image[202];
    assign  image_0_189[55:48]   = Image[203];
    assign  image_0_189[47:40]   = Image[233];
    assign  image_0_189[39:32]   = Image[234];
    assign  image_0_189[31:24]   = Image[235];
    assign  image_0_189[23:16]   = Image[265];
    assign  image_0_189[15:8]    = Image[266];
    assign  image_0_189[7:0]     = Image[267];

    assign  image_0_190[71:64]   = Image[202];
    assign  image_0_190[63:56]   = Image[203];
    assign  image_0_190[55:48]   = Image[204];
    assign  image_0_190[47:40]   = Image[234];
    assign  image_0_190[39:32]   = Image[235];
    assign  image_0_190[31:24]   = Image[236];
    assign  image_0_190[23:16]   = Image[266];
    assign  image_0_190[15:8]    = Image[267];
    assign  image_0_190[7:0]     = Image[268];

    assign  image_0_191[71:64]   = Image[203];
    assign  image_0_191[63:56]   = Image[204];
    assign  image_0_191[55:48]   = Image[205];
    assign  image_0_191[47:40]   = Image[235];
    assign  image_0_191[39:32]   = Image[236];
    assign  image_0_191[31:24]   = Image[237];
    assign  image_0_191[23:16]   = Image[267];
    assign  image_0_191[15:8]    = Image[268];
    assign  image_0_191[7:0]     = Image[269];

    assign  image_0_192[71:64]   = Image[204];
    assign  image_0_192[63:56]   = Image[205];
    assign  image_0_192[55:48]   = Image[206];
    assign  image_0_192[47:40]   = Image[236];
    assign  image_0_192[39:32]   = Image[237];
    assign  image_0_192[31:24]   = Image[238];
    assign  image_0_192[23:16]   = Image[268];
    assign  image_0_192[15:8]    = Image[269];
    assign  image_0_192[7:0]     = Image[270];

    assign  image_0_193[71:64]   = Image[205];
    assign  image_0_193[63:56]   = Image[206];
    assign  image_0_193[55:48]   = Image[207];
    assign  image_0_193[47:40]   = Image[237];
    assign  image_0_193[39:32]   = Image[238];
    assign  image_0_193[31:24]   = Image[239];
    assign  image_0_193[23:16]   = Image[269];
    assign  image_0_193[15:8]    = Image[270];
    assign  image_0_193[7:0]     = Image[271];

    assign  image_0_194[71:64]   = Image[206];
    assign  image_0_194[63:56]   = Image[207];
    assign  image_0_194[55:48]   = Image[208];
    assign  image_0_194[47:40]   = Image[238];
    assign  image_0_194[39:32]   = Image[239];
    assign  image_0_194[31:24]   = Image[240];
    assign  image_0_194[23:16]   = Image[270];
    assign  image_0_194[15:8]    = Image[271];
    assign  image_0_194[7:0]     = Image[272];

    assign  image_0_195[71:64]   = Image[207];
    assign  image_0_195[63:56]   = Image[208];
    assign  image_0_195[55:48]   = Image[209];
    assign  image_0_195[47:40]   = Image[239];
    assign  image_0_195[39:32]   = Image[240];
    assign  image_0_195[31:24]   = Image[241];
    assign  image_0_195[23:16]   = Image[271];
    assign  image_0_195[15:8]    = Image[272];
    assign  image_0_195[7:0]     = Image[273];

    assign  image_0_196[71:64]   = Image[208];
    assign  image_0_196[63:56]   = Image[209];
    assign  image_0_196[55:48]   = Image[210];
    assign  image_0_196[47:40]   = Image[240];
    assign  image_0_196[39:32]   = Image[241];
    assign  image_0_196[31:24]   = Image[242];
    assign  image_0_196[23:16]   = Image[272];
    assign  image_0_196[15:8]    = Image[273];
    assign  image_0_196[7:0]     = Image[274];

    assign  image_0_197[71:64]   = Image[209];
    assign  image_0_197[63:56]   = Image[210];
    assign  image_0_197[55:48]   = Image[211];
    assign  image_0_197[47:40]   = Image[241];
    assign  image_0_197[39:32]   = Image[242];
    assign  image_0_197[31:24]   = Image[243];
    assign  image_0_197[23:16]   = Image[273];
    assign  image_0_197[15:8]    = Image[274];
    assign  image_0_197[7:0]     = Image[275];

    assign  image_0_198[71:64]   = Image[210];
    assign  image_0_198[63:56]   = Image[211];
    assign  image_0_198[55:48]   = Image[212];
    assign  image_0_198[47:40]   = Image[242];
    assign  image_0_198[39:32]   = Image[243];
    assign  image_0_198[31:24]   = Image[244];
    assign  image_0_198[23:16]   = Image[274];
    assign  image_0_198[15:8]    = Image[275];
    assign  image_0_198[7:0]     = Image[276];

    assign  image_0_199[71:64]   = Image[211];
    assign  image_0_199[63:56]   = Image[212];
    assign  image_0_199[55:48]   = Image[213];
    assign  image_0_199[47:40]   = Image[243];
    assign  image_0_199[39:32]   = Image[244];
    assign  image_0_199[31:24]   = Image[245];
    assign  image_0_199[23:16]   = Image[275];
    assign  image_0_199[15:8]    = Image[276];
    assign  image_0_199[7:0]     = Image[277];

    assign  image_0_200[71:64]   = Image[212];
    assign  image_0_200[63:56]   = Image[213];
    assign  image_0_200[55:48]   = Image[214];
    assign  image_0_200[47:40]   = Image[244];
    assign  image_0_200[39:32]   = Image[245];
    assign  image_0_200[31:24]   = Image[246];
    assign  image_0_200[23:16]   = Image[276];
    assign  image_0_200[15:8]    = Image[277];
    assign  image_0_200[7:0]     = Image[278];

    assign  image_0_201[71:64]   = Image[213];
    assign  image_0_201[63:56]   = Image[214];
    assign  image_0_201[55:48]   = Image[215];
    assign  image_0_201[47:40]   = Image[245];
    assign  image_0_201[39:32]   = Image[246];
    assign  image_0_201[31:24]   = Image[247];
    assign  image_0_201[23:16]   = Image[277];
    assign  image_0_201[15:8]    = Image[278];
    assign  image_0_201[7:0]     = Image[279];

    assign  image_0_202[71:64]   = Image[214];
    assign  image_0_202[63:56]   = Image[215];
    assign  image_0_202[55:48]   = Image[216];
    assign  image_0_202[47:40]   = Image[246];
    assign  image_0_202[39:32]   = Image[247];
    assign  image_0_202[31:24]   = Image[248];
    assign  image_0_202[23:16]   = Image[278];
    assign  image_0_202[15:8]    = Image[279];
    assign  image_0_202[7:0]     = Image[280];

    assign  image_0_203[71:64]   = Image[215];
    assign  image_0_203[63:56]   = Image[216];
    assign  image_0_203[55:48]   = Image[217];
    assign  image_0_203[47:40]   = Image[247];
    assign  image_0_203[39:32]   = Image[248];
    assign  image_0_203[31:24]   = Image[249];
    assign  image_0_203[23:16]   = Image[279];
    assign  image_0_203[15:8]    = Image[280];
    assign  image_0_203[7:0]     = Image[281];

    assign  image_0_204[71:64]   = Image[216];
    assign  image_0_204[63:56]   = Image[217];
    assign  image_0_204[55:48]   = Image[218];
    assign  image_0_204[47:40]   = Image[248];
    assign  image_0_204[39:32]   = Image[249];
    assign  image_0_204[31:24]   = Image[250];
    assign  image_0_204[23:16]   = Image[280];
    assign  image_0_204[15:8]    = Image[281];
    assign  image_0_204[7:0]     = Image[282];

    assign  image_0_205[71:64]   = Image[217];
    assign  image_0_205[63:56]   = Image[218];
    assign  image_0_205[55:48]   = Image[219];
    assign  image_0_205[47:40]   = Image[249];
    assign  image_0_205[39:32]   = Image[250];
    assign  image_0_205[31:24]   = Image[251];
    assign  image_0_205[23:16]   = Image[281];
    assign  image_0_205[15:8]    = Image[282];
    assign  image_0_205[7:0]     = Image[283];

    assign  image_0_206[71:64]   = Image[218];
    assign  image_0_206[63:56]   = Image[219];
    assign  image_0_206[55:48]   = Image[220];
    assign  image_0_206[47:40]   = Image[250];
    assign  image_0_206[39:32]   = Image[251];
    assign  image_0_206[31:24]   = Image[252];
    assign  image_0_206[23:16]   = Image[282];
    assign  image_0_206[15:8]    = Image[283];
    assign  image_0_206[7:0]     = Image[284];

    assign  image_0_207[71:64]   = Image[219];
    assign  image_0_207[63:56]   = Image[220];
    assign  image_0_207[55:48]   = Image[221];
    assign  image_0_207[47:40]   = Image[251];
    assign  image_0_207[39:32]   = Image[252];
    assign  image_0_207[31:24]   = Image[253];
    assign  image_0_207[23:16]   = Image[283];
    assign  image_0_207[15:8]    = Image[284];
    assign  image_0_207[7:0]     = Image[285];

    assign  image_0_208[71:64]   = Image[220];
    assign  image_0_208[63:56]   = Image[221];
    assign  image_0_208[55:48]   = Image[222];
    assign  image_0_208[47:40]   = Image[252];
    assign  image_0_208[39:32]   = Image[253];
    assign  image_0_208[31:24]   = Image[254];
    assign  image_0_208[23:16]   = Image[284];
    assign  image_0_208[15:8]    = Image[285];
    assign  image_0_208[7:0]     = Image[286];

    assign  image_0_209[71:64]   = Image[221];
    assign  image_0_209[63:56]   = Image[222];
    assign  image_0_209[55:48]   = Image[223];
    assign  image_0_209[47:40]   = Image[253];
    assign  image_0_209[39:32]   = Image[254];
    assign  image_0_209[31:24]   = Image[255];
    assign  image_0_209[23:16]   = Image[285];
    assign  image_0_209[15:8]    = Image[286];
    assign  image_0_209[7:0]     = Image[287];

    assign  image_0_210[71:64]   = Image[224];
    assign  image_0_210[63:56]   = Image[225];
    assign  image_0_210[55:48]   = Image[226];
    assign  image_0_210[47:40]   = Image[256];
    assign  image_0_210[39:32]   = Image[257];
    assign  image_0_210[31:24]   = Image[258];
    assign  image_0_210[23:16]   = Image[288];
    assign  image_0_210[15:8]    = Image[289];
    assign  image_0_210[7:0]     = Image[290];

    assign  image_0_211[71:64]   = Image[225];
    assign  image_0_211[63:56]   = Image[226];
    assign  image_0_211[55:48]   = Image[227];
    assign  image_0_211[47:40]   = Image[257];
    assign  image_0_211[39:32]   = Image[258];
    assign  image_0_211[31:24]   = Image[259];
    assign  image_0_211[23:16]   = Image[289];
    assign  image_0_211[15:8]    = Image[290];
    assign  image_0_211[7:0]     = Image[291];

    assign  image_0_212[71:64]   = Image[226];
    assign  image_0_212[63:56]   = Image[227];
    assign  image_0_212[55:48]   = Image[228];
    assign  image_0_212[47:40]   = Image[258];
    assign  image_0_212[39:32]   = Image[259];
    assign  image_0_212[31:24]   = Image[260];
    assign  image_0_212[23:16]   = Image[290];
    assign  image_0_212[15:8]    = Image[291];
    assign  image_0_212[7:0]     = Image[292];

    assign  image_0_213[71:64]   = Image[227];
    assign  image_0_213[63:56]   = Image[228];
    assign  image_0_213[55:48]   = Image[229];
    assign  image_0_213[47:40]   = Image[259];
    assign  image_0_213[39:32]   = Image[260];
    assign  image_0_213[31:24]   = Image[261];
    assign  image_0_213[23:16]   = Image[291];
    assign  image_0_213[15:8]    = Image[292];
    assign  image_0_213[7:0]     = Image[293];

    assign  image_0_214[71:64]   = Image[228];
    assign  image_0_214[63:56]   = Image[229];
    assign  image_0_214[55:48]   = Image[230];
    assign  image_0_214[47:40]   = Image[260];
    assign  image_0_214[39:32]   = Image[261];
    assign  image_0_214[31:24]   = Image[262];
    assign  image_0_214[23:16]   = Image[292];
    assign  image_0_214[15:8]    = Image[293];
    assign  image_0_214[7:0]     = Image[294];

    assign  image_0_215[71:64]   = Image[229];
    assign  image_0_215[63:56]   = Image[230];
    assign  image_0_215[55:48]   = Image[231];
    assign  image_0_215[47:40]   = Image[261];
    assign  image_0_215[39:32]   = Image[262];
    assign  image_0_215[31:24]   = Image[263];
    assign  image_0_215[23:16]   = Image[293];
    assign  image_0_215[15:8]    = Image[294];
    assign  image_0_215[7:0]     = Image[295];

    assign  image_0_216[71:64]   = Image[230];
    assign  image_0_216[63:56]   = Image[231];
    assign  image_0_216[55:48]   = Image[232];
    assign  image_0_216[47:40]   = Image[262];
    assign  image_0_216[39:32]   = Image[263];
    assign  image_0_216[31:24]   = Image[264];
    assign  image_0_216[23:16]   = Image[294];
    assign  image_0_216[15:8]    = Image[295];
    assign  image_0_216[7:0]     = Image[296];

    assign  image_0_217[71:64]   = Image[231];
    assign  image_0_217[63:56]   = Image[232];
    assign  image_0_217[55:48]   = Image[233];
    assign  image_0_217[47:40]   = Image[263];
    assign  image_0_217[39:32]   = Image[264];
    assign  image_0_217[31:24]   = Image[265];
    assign  image_0_217[23:16]   = Image[295];
    assign  image_0_217[15:8]    = Image[296];
    assign  image_0_217[7:0]     = Image[297];

    assign  image_0_218[71:64]   = Image[232];
    assign  image_0_218[63:56]   = Image[233];
    assign  image_0_218[55:48]   = Image[234];
    assign  image_0_218[47:40]   = Image[264];
    assign  image_0_218[39:32]   = Image[265];
    assign  image_0_218[31:24]   = Image[266];
    assign  image_0_218[23:16]   = Image[296];
    assign  image_0_218[15:8]    = Image[297];
    assign  image_0_218[7:0]     = Image[298];

    assign  image_0_219[71:64]   = Image[233];
    assign  image_0_219[63:56]   = Image[234];
    assign  image_0_219[55:48]   = Image[235];
    assign  image_0_219[47:40]   = Image[265];
    assign  image_0_219[39:32]   = Image[266];
    assign  image_0_219[31:24]   = Image[267];
    assign  image_0_219[23:16]   = Image[297];
    assign  image_0_219[15:8]    = Image[298];
    assign  image_0_219[7:0]     = Image[299];

    assign  image_0_220[71:64]   = Image[234];
    assign  image_0_220[63:56]   = Image[235];
    assign  image_0_220[55:48]   = Image[236];
    assign  image_0_220[47:40]   = Image[266];
    assign  image_0_220[39:32]   = Image[267];
    assign  image_0_220[31:24]   = Image[268];
    assign  image_0_220[23:16]   = Image[298];
    assign  image_0_220[15:8]    = Image[299];
    assign  image_0_220[7:0]     = Image[300];

    assign  image_0_221[71:64]   = Image[235];
    assign  image_0_221[63:56]   = Image[236];
    assign  image_0_221[55:48]   = Image[237];
    assign  image_0_221[47:40]   = Image[267];
    assign  image_0_221[39:32]   = Image[268];
    assign  image_0_221[31:24]   = Image[269];
    assign  image_0_221[23:16]   = Image[299];
    assign  image_0_221[15:8]    = Image[300];
    assign  image_0_221[7:0]     = Image[301];

    assign  image_0_222[71:64]   = Image[236];
    assign  image_0_222[63:56]   = Image[237];
    assign  image_0_222[55:48]   = Image[238];
    assign  image_0_222[47:40]   = Image[268];
    assign  image_0_222[39:32]   = Image[269];
    assign  image_0_222[31:24]   = Image[270];
    assign  image_0_222[23:16]   = Image[300];
    assign  image_0_222[15:8]    = Image[301];
    assign  image_0_222[7:0]     = Image[302];

    assign  image_0_223[71:64]   = Image[237];
    assign  image_0_223[63:56]   = Image[238];
    assign  image_0_223[55:48]   = Image[239];
    assign  image_0_223[47:40]   = Image[269];
    assign  image_0_223[39:32]   = Image[270];
    assign  image_0_223[31:24]   = Image[271];
    assign  image_0_223[23:16]   = Image[301];
    assign  image_0_223[15:8]    = Image[302];
    assign  image_0_223[7:0]     = Image[303];

    assign  image_0_224[71:64]   = Image[238];
    assign  image_0_224[63:56]   = Image[239];
    assign  image_0_224[55:48]   = Image[240];
    assign  image_0_224[47:40]   = Image[270];
    assign  image_0_224[39:32]   = Image[271];
    assign  image_0_224[31:24]   = Image[272];
    assign  image_0_224[23:16]   = Image[302];
    assign  image_0_224[15:8]    = Image[303];
    assign  image_0_224[7:0]     = Image[304];

    assign  image_0_225[71:64]   = Image[239];
    assign  image_0_225[63:56]   = Image[240];
    assign  image_0_225[55:48]   = Image[241];
    assign  image_0_225[47:40]   = Image[271];
    assign  image_0_225[39:32]   = Image[272];
    assign  image_0_225[31:24]   = Image[273];
    assign  image_0_225[23:16]   = Image[303];
    assign  image_0_225[15:8]    = Image[304];
    assign  image_0_225[7:0]     = Image[305];

    assign  image_0_226[71:64]   = Image[240];
    assign  image_0_226[63:56]   = Image[241];
    assign  image_0_226[55:48]   = Image[242];
    assign  image_0_226[47:40]   = Image[272];
    assign  image_0_226[39:32]   = Image[273];
    assign  image_0_226[31:24]   = Image[274];
    assign  image_0_226[23:16]   = Image[304];
    assign  image_0_226[15:8]    = Image[305];
    assign  image_0_226[7:0]     = Image[306];

    assign  image_0_227[71:64]   = Image[241];
    assign  image_0_227[63:56]   = Image[242];
    assign  image_0_227[55:48]   = Image[243];
    assign  image_0_227[47:40]   = Image[273];
    assign  image_0_227[39:32]   = Image[274];
    assign  image_0_227[31:24]   = Image[275];
    assign  image_0_227[23:16]   = Image[305];
    assign  image_0_227[15:8]    = Image[306];
    assign  image_0_227[7:0]     = Image[307];

    assign  image_0_228[71:64]   = Image[242];
    assign  image_0_228[63:56]   = Image[243];
    assign  image_0_228[55:48]   = Image[244];
    assign  image_0_228[47:40]   = Image[274];
    assign  image_0_228[39:32]   = Image[275];
    assign  image_0_228[31:24]   = Image[276];
    assign  image_0_228[23:16]   = Image[306];
    assign  image_0_228[15:8]    = Image[307];
    assign  image_0_228[7:0]     = Image[308];

    assign  image_0_229[71:64]   = Image[243];
    assign  image_0_229[63:56]   = Image[244];
    assign  image_0_229[55:48]   = Image[245];
    assign  image_0_229[47:40]   = Image[275];
    assign  image_0_229[39:32]   = Image[276];
    assign  image_0_229[31:24]   = Image[277];
    assign  image_0_229[23:16]   = Image[307];
    assign  image_0_229[15:8]    = Image[308];
    assign  image_0_229[7:0]     = Image[309];

    assign  image_0_230[71:64]   = Image[244];
    assign  image_0_230[63:56]   = Image[245];
    assign  image_0_230[55:48]   = Image[246];
    assign  image_0_230[47:40]   = Image[276];
    assign  image_0_230[39:32]   = Image[277];
    assign  image_0_230[31:24]   = Image[278];
    assign  image_0_230[23:16]   = Image[308];
    assign  image_0_230[15:8]    = Image[309];
    assign  image_0_230[7:0]     = Image[310];

    assign  image_0_231[71:64]   = Image[245];
    assign  image_0_231[63:56]   = Image[246];
    assign  image_0_231[55:48]   = Image[247];
    assign  image_0_231[47:40]   = Image[277];
    assign  image_0_231[39:32]   = Image[278];
    assign  image_0_231[31:24]   = Image[279];
    assign  image_0_231[23:16]   = Image[309];
    assign  image_0_231[15:8]    = Image[310];
    assign  image_0_231[7:0]     = Image[311];

    assign  image_0_232[71:64]   = Image[246];
    assign  image_0_232[63:56]   = Image[247];
    assign  image_0_232[55:48]   = Image[248];
    assign  image_0_232[47:40]   = Image[278];
    assign  image_0_232[39:32]   = Image[279];
    assign  image_0_232[31:24]   = Image[280];
    assign  image_0_232[23:16]   = Image[310];
    assign  image_0_232[15:8]    = Image[311];
    assign  image_0_232[7:0]     = Image[312];

    assign  image_0_233[71:64]   = Image[247];
    assign  image_0_233[63:56]   = Image[248];
    assign  image_0_233[55:48]   = Image[249];
    assign  image_0_233[47:40]   = Image[279];
    assign  image_0_233[39:32]   = Image[280];
    assign  image_0_233[31:24]   = Image[281];
    assign  image_0_233[23:16]   = Image[311];
    assign  image_0_233[15:8]    = Image[312];
    assign  image_0_233[7:0]     = Image[313];

    assign  image_0_234[71:64]   = Image[248];
    assign  image_0_234[63:56]   = Image[249];
    assign  image_0_234[55:48]   = Image[250];
    assign  image_0_234[47:40]   = Image[280];
    assign  image_0_234[39:32]   = Image[281];
    assign  image_0_234[31:24]   = Image[282];
    assign  image_0_234[23:16]   = Image[312];
    assign  image_0_234[15:8]    = Image[313];
    assign  image_0_234[7:0]     = Image[314];

    assign  image_0_235[71:64]   = Image[249];
    assign  image_0_235[63:56]   = Image[250];
    assign  image_0_235[55:48]   = Image[251];
    assign  image_0_235[47:40]   = Image[281];
    assign  image_0_235[39:32]   = Image[282];
    assign  image_0_235[31:24]   = Image[283];
    assign  image_0_235[23:16]   = Image[313];
    assign  image_0_235[15:8]    = Image[314];
    assign  image_0_235[7:0]     = Image[315];

    assign  image_0_236[71:64]   = Image[250];
    assign  image_0_236[63:56]   = Image[251];
    assign  image_0_236[55:48]   = Image[252];
    assign  image_0_236[47:40]   = Image[282];
    assign  image_0_236[39:32]   = Image[283];
    assign  image_0_236[31:24]   = Image[284];
    assign  image_0_236[23:16]   = Image[314];
    assign  image_0_236[15:8]    = Image[315];
    assign  image_0_236[7:0]     = Image[316];

    assign  image_0_237[71:64]   = Image[251];
    assign  image_0_237[63:56]   = Image[252];
    assign  image_0_237[55:48]   = Image[253];
    assign  image_0_237[47:40]   = Image[283];
    assign  image_0_237[39:32]   = Image[284];
    assign  image_0_237[31:24]   = Image[285];
    assign  image_0_237[23:16]   = Image[315];
    assign  image_0_237[15:8]    = Image[316];
    assign  image_0_237[7:0]     = Image[317];

    assign  image_0_238[71:64]   = Image[252];
    assign  image_0_238[63:56]   = Image[253];
    assign  image_0_238[55:48]   = Image[254];
    assign  image_0_238[47:40]   = Image[284];
    assign  image_0_238[39:32]   = Image[285];
    assign  image_0_238[31:24]   = Image[286];
    assign  image_0_238[23:16]   = Image[316];
    assign  image_0_238[15:8]    = Image[317];
    assign  image_0_238[7:0]     = Image[318];

    assign  image_0_239[71:64]   = Image[253];
    assign  image_0_239[63:56]   = Image[254];
    assign  image_0_239[55:48]   = Image[255];
    assign  image_0_239[47:40]   = Image[285];
    assign  image_0_239[39:32]   = Image[286];
    assign  image_0_239[31:24]   = Image[287];
    assign  image_0_239[23:16]   = Image[317];
    assign  image_0_239[15:8]    = Image[318];
    assign  image_0_239[7:0]     = Image[319];

    assign  image_0_240[71:64]   = Image[256];
    assign  image_0_240[63:56]   = Image[257];
    assign  image_0_240[55:48]   = Image[258];
    assign  image_0_240[47:40]   = Image[288];
    assign  image_0_240[39:32]   = Image[289];
    assign  image_0_240[31:24]   = Image[290];
    assign  image_0_240[23:16]   = Image[320];
    assign  image_0_240[15:8]    = Image[321];
    assign  image_0_240[7:0]     = Image[322];

    assign  image_0_241[71:64]   = Image[257];
    assign  image_0_241[63:56]   = Image[258];
    assign  image_0_241[55:48]   = Image[259];
    assign  image_0_241[47:40]   = Image[289];
    assign  image_0_241[39:32]   = Image[290];
    assign  image_0_241[31:24]   = Image[291];
    assign  image_0_241[23:16]   = Image[321];
    assign  image_0_241[15:8]    = Image[322];
    assign  image_0_241[7:0]     = Image[323];

    assign  image_0_242[71:64]   = Image[258];
    assign  image_0_242[63:56]   = Image[259];
    assign  image_0_242[55:48]   = Image[260];
    assign  image_0_242[47:40]   = Image[290];
    assign  image_0_242[39:32]   = Image[291];
    assign  image_0_242[31:24]   = Image[292];
    assign  image_0_242[23:16]   = Image[322];
    assign  image_0_242[15:8]    = Image[323];
    assign  image_0_242[7:0]     = Image[324];

    assign  image_0_243[71:64]   = Image[259];
    assign  image_0_243[63:56]   = Image[260];
    assign  image_0_243[55:48]   = Image[261];
    assign  image_0_243[47:40]   = Image[291];
    assign  image_0_243[39:32]   = Image[292];
    assign  image_0_243[31:24]   = Image[293];
    assign  image_0_243[23:16]   = Image[323];
    assign  image_0_243[15:8]    = Image[324];
    assign  image_0_243[7:0]     = Image[325];

    assign  image_0_244[71:64]   = Image[260];
    assign  image_0_244[63:56]   = Image[261];
    assign  image_0_244[55:48]   = Image[262];
    assign  image_0_244[47:40]   = Image[292];
    assign  image_0_244[39:32]   = Image[293];
    assign  image_0_244[31:24]   = Image[294];
    assign  image_0_244[23:16]   = Image[324];
    assign  image_0_244[15:8]    = Image[325];
    assign  image_0_244[7:0]     = Image[326];

    assign  image_0_245[71:64]   = Image[261];
    assign  image_0_245[63:56]   = Image[262];
    assign  image_0_245[55:48]   = Image[263];
    assign  image_0_245[47:40]   = Image[293];
    assign  image_0_245[39:32]   = Image[294];
    assign  image_0_245[31:24]   = Image[295];
    assign  image_0_245[23:16]   = Image[325];
    assign  image_0_245[15:8]    = Image[326];
    assign  image_0_245[7:0]     = Image[327];

    assign  image_0_246[71:64]   = Image[262];
    assign  image_0_246[63:56]   = Image[263];
    assign  image_0_246[55:48]   = Image[264];
    assign  image_0_246[47:40]   = Image[294];
    assign  image_0_246[39:32]   = Image[295];
    assign  image_0_246[31:24]   = Image[296];
    assign  image_0_246[23:16]   = Image[326];
    assign  image_0_246[15:8]    = Image[327];
    assign  image_0_246[7:0]     = Image[328];

    assign  image_0_247[71:64]   = Image[263];
    assign  image_0_247[63:56]   = Image[264];
    assign  image_0_247[55:48]   = Image[265];
    assign  image_0_247[47:40]   = Image[295];
    assign  image_0_247[39:32]   = Image[296];
    assign  image_0_247[31:24]   = Image[297];
    assign  image_0_247[23:16]   = Image[327];
    assign  image_0_247[15:8]    = Image[328];
    assign  image_0_247[7:0]     = Image[329];

    assign  image_0_248[71:64]   = Image[264];
    assign  image_0_248[63:56]   = Image[265];
    assign  image_0_248[55:48]   = Image[266];
    assign  image_0_248[47:40]   = Image[296];
    assign  image_0_248[39:32]   = Image[297];
    assign  image_0_248[31:24]   = Image[298];
    assign  image_0_248[23:16]   = Image[328];
    assign  image_0_248[15:8]    = Image[329];
    assign  image_0_248[7:0]     = Image[330];

    assign  image_0_249[71:64]   = Image[265];
    assign  image_0_249[63:56]   = Image[266];
    assign  image_0_249[55:48]   = Image[267];
    assign  image_0_249[47:40]   = Image[297];
    assign  image_0_249[39:32]   = Image[298];
    assign  image_0_249[31:24]   = Image[299];
    assign  image_0_249[23:16]   = Image[329];
    assign  image_0_249[15:8]    = Image[330];
    assign  image_0_249[7:0]     = Image[331];

    assign  image_0_250[71:64]   = Image[266];
    assign  image_0_250[63:56]   = Image[267];
    assign  image_0_250[55:48]   = Image[268];
    assign  image_0_250[47:40]   = Image[298];
    assign  image_0_250[39:32]   = Image[299];
    assign  image_0_250[31:24]   = Image[300];
    assign  image_0_250[23:16]   = Image[330];
    assign  image_0_250[15:8]    = Image[331];
    assign  image_0_250[7:0]     = Image[332];

    assign  image_0_251[71:64]   = Image[267];
    assign  image_0_251[63:56]   = Image[268];
    assign  image_0_251[55:48]   = Image[269];
    assign  image_0_251[47:40]   = Image[299];
    assign  image_0_251[39:32]   = Image[300];
    assign  image_0_251[31:24]   = Image[301];
    assign  image_0_251[23:16]   = Image[331];
    assign  image_0_251[15:8]    = Image[332];
    assign  image_0_251[7:0]     = Image[333];

    assign  image_0_252[71:64]   = Image[268];
    assign  image_0_252[63:56]   = Image[269];
    assign  image_0_252[55:48]   = Image[270];
    assign  image_0_252[47:40]   = Image[300];
    assign  image_0_252[39:32]   = Image[301];
    assign  image_0_252[31:24]   = Image[302];
    assign  image_0_252[23:16]   = Image[332];
    assign  image_0_252[15:8]    = Image[333];
    assign  image_0_252[7:0]     = Image[334];

    assign  image_0_253[71:64]   = Image[269];
    assign  image_0_253[63:56]   = Image[270];
    assign  image_0_253[55:48]   = Image[271];
    assign  image_0_253[47:40]   = Image[301];
    assign  image_0_253[39:32]   = Image[302];
    assign  image_0_253[31:24]   = Image[303];
    assign  image_0_253[23:16]   = Image[333];
    assign  image_0_253[15:8]    = Image[334];
    assign  image_0_253[7:0]     = Image[335];

    assign  image_0_254[71:64]   = Image[270];
    assign  image_0_254[63:56]   = Image[271];
    assign  image_0_254[55:48]   = Image[272];
    assign  image_0_254[47:40]   = Image[302];
    assign  image_0_254[39:32]   = Image[303];
    assign  image_0_254[31:24]   = Image[304];
    assign  image_0_254[23:16]   = Image[334];
    assign  image_0_254[15:8]    = Image[335];
    assign  image_0_254[7:0]     = Image[336];

    assign  image_0_255[71:64]   = Image[271];
    assign  image_0_255[63:56]   = Image[272];
    assign  image_0_255[55:48]   = Image[273];
    assign  image_0_255[47:40]   = Image[303];
    assign  image_0_255[39:32]   = Image[304];
    assign  image_0_255[31:24]   = Image[305];
    assign  image_0_255[23:16]   = Image[335];
    assign  image_0_255[15:8]    = Image[336];
    assign  image_0_255[7:0]     = Image[337];

    assign  image_0_256[71:64]   = Image[272];
    assign  image_0_256[63:56]   = Image[273];
    assign  image_0_256[55:48]   = Image[274];
    assign  image_0_256[47:40]   = Image[304];
    assign  image_0_256[39:32]   = Image[305];
    assign  image_0_256[31:24]   = Image[306];
    assign  image_0_256[23:16]   = Image[336];
    assign  image_0_256[15:8]    = Image[337];
    assign  image_0_256[7:0]     = Image[338];

    assign  image_0_257[71:64]   = Image[273];
    assign  image_0_257[63:56]   = Image[274];
    assign  image_0_257[55:48]   = Image[275];
    assign  image_0_257[47:40]   = Image[305];
    assign  image_0_257[39:32]   = Image[306];
    assign  image_0_257[31:24]   = Image[307];
    assign  image_0_257[23:16]   = Image[337];
    assign  image_0_257[15:8]    = Image[338];
    assign  image_0_257[7:0]     = Image[339];

    assign  image_0_258[71:64]   = Image[274];
    assign  image_0_258[63:56]   = Image[275];
    assign  image_0_258[55:48]   = Image[276];
    assign  image_0_258[47:40]   = Image[306];
    assign  image_0_258[39:32]   = Image[307];
    assign  image_0_258[31:24]   = Image[308];
    assign  image_0_258[23:16]   = Image[338];
    assign  image_0_258[15:8]    = Image[339];
    assign  image_0_258[7:0]     = Image[340];

    assign  image_0_259[71:64]   = Image[275];
    assign  image_0_259[63:56]   = Image[276];
    assign  image_0_259[55:48]   = Image[277];
    assign  image_0_259[47:40]   = Image[307];
    assign  image_0_259[39:32]   = Image[308];
    assign  image_0_259[31:24]   = Image[309];
    assign  image_0_259[23:16]   = Image[339];
    assign  image_0_259[15:8]    = Image[340];
    assign  image_0_259[7:0]     = Image[341];

    assign  image_0_260[71:64]   = Image[276];
    assign  image_0_260[63:56]   = Image[277];
    assign  image_0_260[55:48]   = Image[278];
    assign  image_0_260[47:40]   = Image[308];
    assign  image_0_260[39:32]   = Image[309];
    assign  image_0_260[31:24]   = Image[310];
    assign  image_0_260[23:16]   = Image[340];
    assign  image_0_260[15:8]    = Image[341];
    assign  image_0_260[7:0]     = Image[342];

    assign  image_0_261[71:64]   = Image[277];
    assign  image_0_261[63:56]   = Image[278];
    assign  image_0_261[55:48]   = Image[279];
    assign  image_0_261[47:40]   = Image[309];
    assign  image_0_261[39:32]   = Image[310];
    assign  image_0_261[31:24]   = Image[311];
    assign  image_0_261[23:16]   = Image[341];
    assign  image_0_261[15:8]    = Image[342];
    assign  image_0_261[7:0]     = Image[343];

    assign  image_0_262[71:64]   = Image[278];
    assign  image_0_262[63:56]   = Image[279];
    assign  image_0_262[55:48]   = Image[280];
    assign  image_0_262[47:40]   = Image[310];
    assign  image_0_262[39:32]   = Image[311];
    assign  image_0_262[31:24]   = Image[312];
    assign  image_0_262[23:16]   = Image[342];
    assign  image_0_262[15:8]    = Image[343];
    assign  image_0_262[7:0]     = Image[344];

    assign  image_0_263[71:64]   = Image[279];
    assign  image_0_263[63:56]   = Image[280];
    assign  image_0_263[55:48]   = Image[281];
    assign  image_0_263[47:40]   = Image[311];
    assign  image_0_263[39:32]   = Image[312];
    assign  image_0_263[31:24]   = Image[313];
    assign  image_0_263[23:16]   = Image[343];
    assign  image_0_263[15:8]    = Image[344];
    assign  image_0_263[7:0]     = Image[345];

    assign  image_0_264[71:64]   = Image[280];
    assign  image_0_264[63:56]   = Image[281];
    assign  image_0_264[55:48]   = Image[282];
    assign  image_0_264[47:40]   = Image[312];
    assign  image_0_264[39:32]   = Image[313];
    assign  image_0_264[31:24]   = Image[314];
    assign  image_0_264[23:16]   = Image[344];
    assign  image_0_264[15:8]    = Image[345];
    assign  image_0_264[7:0]     = Image[346];

    assign  image_0_265[71:64]   = Image[281];
    assign  image_0_265[63:56]   = Image[282];
    assign  image_0_265[55:48]   = Image[283];
    assign  image_0_265[47:40]   = Image[313];
    assign  image_0_265[39:32]   = Image[314];
    assign  image_0_265[31:24]   = Image[315];
    assign  image_0_265[23:16]   = Image[345];
    assign  image_0_265[15:8]    = Image[346];
    assign  image_0_265[7:0]     = Image[347];

    assign  image_0_266[71:64]   = Image[282];
    assign  image_0_266[63:56]   = Image[283];
    assign  image_0_266[55:48]   = Image[284];
    assign  image_0_266[47:40]   = Image[314];
    assign  image_0_266[39:32]   = Image[315];
    assign  image_0_266[31:24]   = Image[316];
    assign  image_0_266[23:16]   = Image[346];
    assign  image_0_266[15:8]    = Image[347];
    assign  image_0_266[7:0]     = Image[348];

    assign  image_0_267[71:64]   = Image[283];
    assign  image_0_267[63:56]   = Image[284];
    assign  image_0_267[55:48]   = Image[285];
    assign  image_0_267[47:40]   = Image[315];
    assign  image_0_267[39:32]   = Image[316];
    assign  image_0_267[31:24]   = Image[317];
    assign  image_0_267[23:16]   = Image[347];
    assign  image_0_267[15:8]    = Image[348];
    assign  image_0_267[7:0]     = Image[349];

    assign  image_0_268[71:64]   = Image[284];
    assign  image_0_268[63:56]   = Image[285];
    assign  image_0_268[55:48]   = Image[286];
    assign  image_0_268[47:40]   = Image[316];
    assign  image_0_268[39:32]   = Image[317];
    assign  image_0_268[31:24]   = Image[318];
    assign  image_0_268[23:16]   = Image[348];
    assign  image_0_268[15:8]    = Image[349];
    assign  image_0_268[7:0]     = Image[350];

    assign  image_0_269[71:64]   = Image[285];
    assign  image_0_269[63:56]   = Image[286];
    assign  image_0_269[55:48]   = Image[287];
    assign  image_0_269[47:40]   = Image[317];
    assign  image_0_269[39:32]   = Image[318];
    assign  image_0_269[31:24]   = Image[319];
    assign  image_0_269[23:16]   = Image[349];
    assign  image_0_269[15:8]    = Image[350];
    assign  image_0_269[7:0]     = Image[351];

    assign  image_0_270[71:64]   = Image[288];
    assign  image_0_270[63:56]   = Image[289];
    assign  image_0_270[55:48]   = Image[290];
    assign  image_0_270[47:40]   = Image[320];
    assign  image_0_270[39:32]   = Image[321];
    assign  image_0_270[31:24]   = Image[322];
    assign  image_0_270[23:16]   = Image[352];
    assign  image_0_270[15:8]    = Image[353];
    assign  image_0_270[7:0]     = Image[354];

    assign  image_0_271[71:64]   = Image[289];
    assign  image_0_271[63:56]   = Image[290];
    assign  image_0_271[55:48]   = Image[291];
    assign  image_0_271[47:40]   = Image[321];
    assign  image_0_271[39:32]   = Image[322];
    assign  image_0_271[31:24]   = Image[323];
    assign  image_0_271[23:16]   = Image[353];
    assign  image_0_271[15:8]    = Image[354];
    assign  image_0_271[7:0]     = Image[355];

    assign  image_0_272[71:64]   = Image[290];
    assign  image_0_272[63:56]   = Image[291];
    assign  image_0_272[55:48]   = Image[292];
    assign  image_0_272[47:40]   = Image[322];
    assign  image_0_272[39:32]   = Image[323];
    assign  image_0_272[31:24]   = Image[324];
    assign  image_0_272[23:16]   = Image[354];
    assign  image_0_272[15:8]    = Image[355];
    assign  image_0_272[7:0]     = Image[356];

    assign  image_0_273[71:64]   = Image[291];
    assign  image_0_273[63:56]   = Image[292];
    assign  image_0_273[55:48]   = Image[293];
    assign  image_0_273[47:40]   = Image[323];
    assign  image_0_273[39:32]   = Image[324];
    assign  image_0_273[31:24]   = Image[325];
    assign  image_0_273[23:16]   = Image[355];
    assign  image_0_273[15:8]    = Image[356];
    assign  image_0_273[7:0]     = Image[357];

    assign  image_0_274[71:64]   = Image[292];
    assign  image_0_274[63:56]   = Image[293];
    assign  image_0_274[55:48]   = Image[294];
    assign  image_0_274[47:40]   = Image[324];
    assign  image_0_274[39:32]   = Image[325];
    assign  image_0_274[31:24]   = Image[326];
    assign  image_0_274[23:16]   = Image[356];
    assign  image_0_274[15:8]    = Image[357];
    assign  image_0_274[7:0]     = Image[358];

    assign  image_0_275[71:64]   = Image[293];
    assign  image_0_275[63:56]   = Image[294];
    assign  image_0_275[55:48]   = Image[295];
    assign  image_0_275[47:40]   = Image[325];
    assign  image_0_275[39:32]   = Image[326];
    assign  image_0_275[31:24]   = Image[327];
    assign  image_0_275[23:16]   = Image[357];
    assign  image_0_275[15:8]    = Image[358];
    assign  image_0_275[7:0]     = Image[359];

    assign  image_0_276[71:64]   = Image[294];
    assign  image_0_276[63:56]   = Image[295];
    assign  image_0_276[55:48]   = Image[296];
    assign  image_0_276[47:40]   = Image[326];
    assign  image_0_276[39:32]   = Image[327];
    assign  image_0_276[31:24]   = Image[328];
    assign  image_0_276[23:16]   = Image[358];
    assign  image_0_276[15:8]    = Image[359];
    assign  image_0_276[7:0]     = Image[360];

    assign  image_0_277[71:64]   = Image[295];
    assign  image_0_277[63:56]   = Image[296];
    assign  image_0_277[55:48]   = Image[297];
    assign  image_0_277[47:40]   = Image[327];
    assign  image_0_277[39:32]   = Image[328];
    assign  image_0_277[31:24]   = Image[329];
    assign  image_0_277[23:16]   = Image[359];
    assign  image_0_277[15:8]    = Image[360];
    assign  image_0_277[7:0]     = Image[361];

    assign  image_0_278[71:64]   = Image[296];
    assign  image_0_278[63:56]   = Image[297];
    assign  image_0_278[55:48]   = Image[298];
    assign  image_0_278[47:40]   = Image[328];
    assign  image_0_278[39:32]   = Image[329];
    assign  image_0_278[31:24]   = Image[330];
    assign  image_0_278[23:16]   = Image[360];
    assign  image_0_278[15:8]    = Image[361];
    assign  image_0_278[7:0]     = Image[362];

    assign  image_0_279[71:64]   = Image[297];
    assign  image_0_279[63:56]   = Image[298];
    assign  image_0_279[55:48]   = Image[299];
    assign  image_0_279[47:40]   = Image[329];
    assign  image_0_279[39:32]   = Image[330];
    assign  image_0_279[31:24]   = Image[331];
    assign  image_0_279[23:16]   = Image[361];
    assign  image_0_279[15:8]    = Image[362];
    assign  image_0_279[7:0]     = Image[363];

    assign  image_0_280[71:64]   = Image[298];
    assign  image_0_280[63:56]   = Image[299];
    assign  image_0_280[55:48]   = Image[300];
    assign  image_0_280[47:40]   = Image[330];
    assign  image_0_280[39:32]   = Image[331];
    assign  image_0_280[31:24]   = Image[332];
    assign  image_0_280[23:16]   = Image[362];
    assign  image_0_280[15:8]    = Image[363];
    assign  image_0_280[7:0]     = Image[364];

    assign  image_0_281[71:64]   = Image[299];
    assign  image_0_281[63:56]   = Image[300];
    assign  image_0_281[55:48]   = Image[301];
    assign  image_0_281[47:40]   = Image[331];
    assign  image_0_281[39:32]   = Image[332];
    assign  image_0_281[31:24]   = Image[333];
    assign  image_0_281[23:16]   = Image[363];
    assign  image_0_281[15:8]    = Image[364];
    assign  image_0_281[7:0]     = Image[365];

    assign  image_0_282[71:64]   = Image[300];
    assign  image_0_282[63:56]   = Image[301];
    assign  image_0_282[55:48]   = Image[302];
    assign  image_0_282[47:40]   = Image[332];
    assign  image_0_282[39:32]   = Image[333];
    assign  image_0_282[31:24]   = Image[334];
    assign  image_0_282[23:16]   = Image[364];
    assign  image_0_282[15:8]    = Image[365];
    assign  image_0_282[7:0]     = Image[366];

    assign  image_0_283[71:64]   = Image[301];
    assign  image_0_283[63:56]   = Image[302];
    assign  image_0_283[55:48]   = Image[303];
    assign  image_0_283[47:40]   = Image[333];
    assign  image_0_283[39:32]   = Image[334];
    assign  image_0_283[31:24]   = Image[335];
    assign  image_0_283[23:16]   = Image[365];
    assign  image_0_283[15:8]    = Image[366];
    assign  image_0_283[7:0]     = Image[367];

    assign  image_0_284[71:64]   = Image[302];
    assign  image_0_284[63:56]   = Image[303];
    assign  image_0_284[55:48]   = Image[304];
    assign  image_0_284[47:40]   = Image[334];
    assign  image_0_284[39:32]   = Image[335];
    assign  image_0_284[31:24]   = Image[336];
    assign  image_0_284[23:16]   = Image[366];
    assign  image_0_284[15:8]    = Image[367];
    assign  image_0_284[7:0]     = Image[368];

    assign  image_0_285[71:64]   = Image[303];
    assign  image_0_285[63:56]   = Image[304];
    assign  image_0_285[55:48]   = Image[305];
    assign  image_0_285[47:40]   = Image[335];
    assign  image_0_285[39:32]   = Image[336];
    assign  image_0_285[31:24]   = Image[337];
    assign  image_0_285[23:16]   = Image[367];
    assign  image_0_285[15:8]    = Image[368];
    assign  image_0_285[7:0]     = Image[369];

    assign  image_0_286[71:64]   = Image[304];
    assign  image_0_286[63:56]   = Image[305];
    assign  image_0_286[55:48]   = Image[306];
    assign  image_0_286[47:40]   = Image[336];
    assign  image_0_286[39:32]   = Image[337];
    assign  image_0_286[31:24]   = Image[338];
    assign  image_0_286[23:16]   = Image[368];
    assign  image_0_286[15:8]    = Image[369];
    assign  image_0_286[7:0]     = Image[370];

    assign  image_0_287[71:64]   = Image[305];
    assign  image_0_287[63:56]   = Image[306];
    assign  image_0_287[55:48]   = Image[307];
    assign  image_0_287[47:40]   = Image[337];
    assign  image_0_287[39:32]   = Image[338];
    assign  image_0_287[31:24]   = Image[339];
    assign  image_0_287[23:16]   = Image[369];
    assign  image_0_287[15:8]    = Image[370];
    assign  image_0_287[7:0]     = Image[371];

    assign  image_0_288[71:64]   = Image[306];
    assign  image_0_288[63:56]   = Image[307];
    assign  image_0_288[55:48]   = Image[308];
    assign  image_0_288[47:40]   = Image[338];
    assign  image_0_288[39:32]   = Image[339];
    assign  image_0_288[31:24]   = Image[340];
    assign  image_0_288[23:16]   = Image[370];
    assign  image_0_288[15:8]    = Image[371];
    assign  image_0_288[7:0]     = Image[372];

    assign  image_0_289[71:64]   = Image[307];
    assign  image_0_289[63:56]   = Image[308];
    assign  image_0_289[55:48]   = Image[309];
    assign  image_0_289[47:40]   = Image[339];
    assign  image_0_289[39:32]   = Image[340];
    assign  image_0_289[31:24]   = Image[341];
    assign  image_0_289[23:16]   = Image[371];
    assign  image_0_289[15:8]    = Image[372];
    assign  image_0_289[7:0]     = Image[373];

    assign  image_0_290[71:64]   = Image[308];
    assign  image_0_290[63:56]   = Image[309];
    assign  image_0_290[55:48]   = Image[310];
    assign  image_0_290[47:40]   = Image[340];
    assign  image_0_290[39:32]   = Image[341];
    assign  image_0_290[31:24]   = Image[342];
    assign  image_0_290[23:16]   = Image[372];
    assign  image_0_290[15:8]    = Image[373];
    assign  image_0_290[7:0]     = Image[374];

    assign  image_0_291[71:64]   = Image[309];
    assign  image_0_291[63:56]   = Image[310];
    assign  image_0_291[55:48]   = Image[311];
    assign  image_0_291[47:40]   = Image[341];
    assign  image_0_291[39:32]   = Image[342];
    assign  image_0_291[31:24]   = Image[343];
    assign  image_0_291[23:16]   = Image[373];
    assign  image_0_291[15:8]    = Image[374];
    assign  image_0_291[7:0]     = Image[375];

    assign  image_0_292[71:64]   = Image[310];
    assign  image_0_292[63:56]   = Image[311];
    assign  image_0_292[55:48]   = Image[312];
    assign  image_0_292[47:40]   = Image[342];
    assign  image_0_292[39:32]   = Image[343];
    assign  image_0_292[31:24]   = Image[344];
    assign  image_0_292[23:16]   = Image[374];
    assign  image_0_292[15:8]    = Image[375];
    assign  image_0_292[7:0]     = Image[376];

    assign  image_0_293[71:64]   = Image[311];
    assign  image_0_293[63:56]   = Image[312];
    assign  image_0_293[55:48]   = Image[313];
    assign  image_0_293[47:40]   = Image[343];
    assign  image_0_293[39:32]   = Image[344];
    assign  image_0_293[31:24]   = Image[345];
    assign  image_0_293[23:16]   = Image[375];
    assign  image_0_293[15:8]    = Image[376];
    assign  image_0_293[7:0]     = Image[377];

    assign  image_0_294[71:64]   = Image[312];
    assign  image_0_294[63:56]   = Image[313];
    assign  image_0_294[55:48]   = Image[314];
    assign  image_0_294[47:40]   = Image[344];
    assign  image_0_294[39:32]   = Image[345];
    assign  image_0_294[31:24]   = Image[346];
    assign  image_0_294[23:16]   = Image[376];
    assign  image_0_294[15:8]    = Image[377];
    assign  image_0_294[7:0]     = Image[378];

    assign  image_0_295[71:64]   = Image[313];
    assign  image_0_295[63:56]   = Image[314];
    assign  image_0_295[55:48]   = Image[315];
    assign  image_0_295[47:40]   = Image[345];
    assign  image_0_295[39:32]   = Image[346];
    assign  image_0_295[31:24]   = Image[347];
    assign  image_0_295[23:16]   = Image[377];
    assign  image_0_295[15:8]    = Image[378];
    assign  image_0_295[7:0]     = Image[379];

    assign  image_0_296[71:64]   = Image[314];
    assign  image_0_296[63:56]   = Image[315];
    assign  image_0_296[55:48]   = Image[316];
    assign  image_0_296[47:40]   = Image[346];
    assign  image_0_296[39:32]   = Image[347];
    assign  image_0_296[31:24]   = Image[348];
    assign  image_0_296[23:16]   = Image[378];
    assign  image_0_296[15:8]    = Image[379];
    assign  image_0_296[7:0]     = Image[380];

    assign  image_0_297[71:64]   = Image[315];
    assign  image_0_297[63:56]   = Image[316];
    assign  image_0_297[55:48]   = Image[317];
    assign  image_0_297[47:40]   = Image[347];
    assign  image_0_297[39:32]   = Image[348];
    assign  image_0_297[31:24]   = Image[349];
    assign  image_0_297[23:16]   = Image[379];
    assign  image_0_297[15:8]    = Image[380];
    assign  image_0_297[7:0]     = Image[381];

    assign  image_0_298[71:64]   = Image[316];
    assign  image_0_298[63:56]   = Image[317];
    assign  image_0_298[55:48]   = Image[318];
    assign  image_0_298[47:40]   = Image[348];
    assign  image_0_298[39:32]   = Image[349];
    assign  image_0_298[31:24]   = Image[350];
    assign  image_0_298[23:16]   = Image[380];
    assign  image_0_298[15:8]    = Image[381];
    assign  image_0_298[7:0]     = Image[382];

    assign  image_0_299[71:64]   = Image[317];
    assign  image_0_299[63:56]   = Image[318];
    assign  image_0_299[55:48]   = Image[319];
    assign  image_0_299[47:40]   = Image[349];
    assign  image_0_299[39:32]   = Image[350];
    assign  image_0_299[31:24]   = Image[351];
    assign  image_0_299[23:16]   = Image[381];
    assign  image_0_299[15:8]    = Image[382];
    assign  image_0_299[7:0]     = Image[383];

    assign  image_0_300[71:64]   = Image[320];
    assign  image_0_300[63:56]   = Image[321];
    assign  image_0_300[55:48]   = Image[322];
    assign  image_0_300[47:40]   = Image[352];
    assign  image_0_300[39:32]   = Image[353];
    assign  image_0_300[31:24]   = Image[354];
    assign  image_0_300[23:16]   = Image[384];
    assign  image_0_300[15:8]    = Image[385];
    assign  image_0_300[7:0]     = Image[386];

    assign  image_0_301[71:64]   = Image[321];
    assign  image_0_301[63:56]   = Image[322];
    assign  image_0_301[55:48]   = Image[323];
    assign  image_0_301[47:40]   = Image[353];
    assign  image_0_301[39:32]   = Image[354];
    assign  image_0_301[31:24]   = Image[355];
    assign  image_0_301[23:16]   = Image[385];
    assign  image_0_301[15:8]    = Image[386];
    assign  image_0_301[7:0]     = Image[387];

    assign  image_0_302[71:64]   = Image[322];
    assign  image_0_302[63:56]   = Image[323];
    assign  image_0_302[55:48]   = Image[324];
    assign  image_0_302[47:40]   = Image[354];
    assign  image_0_302[39:32]   = Image[355];
    assign  image_0_302[31:24]   = Image[356];
    assign  image_0_302[23:16]   = Image[386];
    assign  image_0_302[15:8]    = Image[387];
    assign  image_0_302[7:0]     = Image[388];

    assign  image_0_303[71:64]   = Image[323];
    assign  image_0_303[63:56]   = Image[324];
    assign  image_0_303[55:48]   = Image[325];
    assign  image_0_303[47:40]   = Image[355];
    assign  image_0_303[39:32]   = Image[356];
    assign  image_0_303[31:24]   = Image[357];
    assign  image_0_303[23:16]   = Image[387];
    assign  image_0_303[15:8]    = Image[388];
    assign  image_0_303[7:0]     = Image[389];

    assign  image_0_304[71:64]   = Image[324];
    assign  image_0_304[63:56]   = Image[325];
    assign  image_0_304[55:48]   = Image[326];
    assign  image_0_304[47:40]   = Image[356];
    assign  image_0_304[39:32]   = Image[357];
    assign  image_0_304[31:24]   = Image[358];
    assign  image_0_304[23:16]   = Image[388];
    assign  image_0_304[15:8]    = Image[389];
    assign  image_0_304[7:0]     = Image[390];

    assign  image_0_305[71:64]   = Image[325];
    assign  image_0_305[63:56]   = Image[326];
    assign  image_0_305[55:48]   = Image[327];
    assign  image_0_305[47:40]   = Image[357];
    assign  image_0_305[39:32]   = Image[358];
    assign  image_0_305[31:24]   = Image[359];
    assign  image_0_305[23:16]   = Image[389];
    assign  image_0_305[15:8]    = Image[390];
    assign  image_0_305[7:0]     = Image[391];

    assign  image_0_306[71:64]   = Image[326];
    assign  image_0_306[63:56]   = Image[327];
    assign  image_0_306[55:48]   = Image[328];
    assign  image_0_306[47:40]   = Image[358];
    assign  image_0_306[39:32]   = Image[359];
    assign  image_0_306[31:24]   = Image[360];
    assign  image_0_306[23:16]   = Image[390];
    assign  image_0_306[15:8]    = Image[391];
    assign  image_0_306[7:0]     = Image[392];

    assign  image_0_307[71:64]   = Image[327];
    assign  image_0_307[63:56]   = Image[328];
    assign  image_0_307[55:48]   = Image[329];
    assign  image_0_307[47:40]   = Image[359];
    assign  image_0_307[39:32]   = Image[360];
    assign  image_0_307[31:24]   = Image[361];
    assign  image_0_307[23:16]   = Image[391];
    assign  image_0_307[15:8]    = Image[392];
    assign  image_0_307[7:0]     = Image[393];

    assign  image_0_308[71:64]   = Image[328];
    assign  image_0_308[63:56]   = Image[329];
    assign  image_0_308[55:48]   = Image[330];
    assign  image_0_308[47:40]   = Image[360];
    assign  image_0_308[39:32]   = Image[361];
    assign  image_0_308[31:24]   = Image[362];
    assign  image_0_308[23:16]   = Image[392];
    assign  image_0_308[15:8]    = Image[393];
    assign  image_0_308[7:0]     = Image[394];

    assign  image_0_309[71:64]   = Image[329];
    assign  image_0_309[63:56]   = Image[330];
    assign  image_0_309[55:48]   = Image[331];
    assign  image_0_309[47:40]   = Image[361];
    assign  image_0_309[39:32]   = Image[362];
    assign  image_0_309[31:24]   = Image[363];
    assign  image_0_309[23:16]   = Image[393];
    assign  image_0_309[15:8]    = Image[394];
    assign  image_0_309[7:0]     = Image[395];

    assign  image_0_310[71:64]   = Image[330];
    assign  image_0_310[63:56]   = Image[331];
    assign  image_0_310[55:48]   = Image[332];
    assign  image_0_310[47:40]   = Image[362];
    assign  image_0_310[39:32]   = Image[363];
    assign  image_0_310[31:24]   = Image[364];
    assign  image_0_310[23:16]   = Image[394];
    assign  image_0_310[15:8]    = Image[395];
    assign  image_0_310[7:0]     = Image[396];

    assign  image_0_311[71:64]   = Image[331];
    assign  image_0_311[63:56]   = Image[332];
    assign  image_0_311[55:48]   = Image[333];
    assign  image_0_311[47:40]   = Image[363];
    assign  image_0_311[39:32]   = Image[364];
    assign  image_0_311[31:24]   = Image[365];
    assign  image_0_311[23:16]   = Image[395];
    assign  image_0_311[15:8]    = Image[396];
    assign  image_0_311[7:0]     = Image[397];

    assign  image_0_312[71:64]   = Image[332];
    assign  image_0_312[63:56]   = Image[333];
    assign  image_0_312[55:48]   = Image[334];
    assign  image_0_312[47:40]   = Image[364];
    assign  image_0_312[39:32]   = Image[365];
    assign  image_0_312[31:24]   = Image[366];
    assign  image_0_312[23:16]   = Image[396];
    assign  image_0_312[15:8]    = Image[397];
    assign  image_0_312[7:0]     = Image[398];

    assign  image_0_313[71:64]   = Image[333];
    assign  image_0_313[63:56]   = Image[334];
    assign  image_0_313[55:48]   = Image[335];
    assign  image_0_313[47:40]   = Image[365];
    assign  image_0_313[39:32]   = Image[366];
    assign  image_0_313[31:24]   = Image[367];
    assign  image_0_313[23:16]   = Image[397];
    assign  image_0_313[15:8]    = Image[398];
    assign  image_0_313[7:0]     = Image[399];

    assign  image_0_314[71:64]   = Image[334];
    assign  image_0_314[63:56]   = Image[335];
    assign  image_0_314[55:48]   = Image[336];
    assign  image_0_314[47:40]   = Image[366];
    assign  image_0_314[39:32]   = Image[367];
    assign  image_0_314[31:24]   = Image[368];
    assign  image_0_314[23:16]   = Image[398];
    assign  image_0_314[15:8]    = Image[399];
    assign  image_0_314[7:0]     = Image[400];

    assign  image_0_315[71:64]   = Image[335];
    assign  image_0_315[63:56]   = Image[336];
    assign  image_0_315[55:48]   = Image[337];
    assign  image_0_315[47:40]   = Image[367];
    assign  image_0_315[39:32]   = Image[368];
    assign  image_0_315[31:24]   = Image[369];
    assign  image_0_315[23:16]   = Image[399];
    assign  image_0_315[15:8]    = Image[400];
    assign  image_0_315[7:0]     = Image[401];

    assign  image_0_316[71:64]   = Image[336];
    assign  image_0_316[63:56]   = Image[337];
    assign  image_0_316[55:48]   = Image[338];
    assign  image_0_316[47:40]   = Image[368];
    assign  image_0_316[39:32]   = Image[369];
    assign  image_0_316[31:24]   = Image[370];
    assign  image_0_316[23:16]   = Image[400];
    assign  image_0_316[15:8]    = Image[401];
    assign  image_0_316[7:0]     = Image[402];

    assign  image_0_317[71:64]   = Image[337];
    assign  image_0_317[63:56]   = Image[338];
    assign  image_0_317[55:48]   = Image[339];
    assign  image_0_317[47:40]   = Image[369];
    assign  image_0_317[39:32]   = Image[370];
    assign  image_0_317[31:24]   = Image[371];
    assign  image_0_317[23:16]   = Image[401];
    assign  image_0_317[15:8]    = Image[402];
    assign  image_0_317[7:0]     = Image[403];

    assign  image_0_318[71:64]   = Image[338];
    assign  image_0_318[63:56]   = Image[339];
    assign  image_0_318[55:48]   = Image[340];
    assign  image_0_318[47:40]   = Image[370];
    assign  image_0_318[39:32]   = Image[371];
    assign  image_0_318[31:24]   = Image[372];
    assign  image_0_318[23:16]   = Image[402];
    assign  image_0_318[15:8]    = Image[403];
    assign  image_0_318[7:0]     = Image[404];

    assign  image_0_319[71:64]   = Image[339];
    assign  image_0_319[63:56]   = Image[340];
    assign  image_0_319[55:48]   = Image[341];
    assign  image_0_319[47:40]   = Image[371];
    assign  image_0_319[39:32]   = Image[372];
    assign  image_0_319[31:24]   = Image[373];
    assign  image_0_319[23:16]   = Image[403];
    assign  image_0_319[15:8]    = Image[404];
    assign  image_0_319[7:0]     = Image[405];

    assign  image_0_320[71:64]   = Image[340];
    assign  image_0_320[63:56]   = Image[341];
    assign  image_0_320[55:48]   = Image[342];
    assign  image_0_320[47:40]   = Image[372];
    assign  image_0_320[39:32]   = Image[373];
    assign  image_0_320[31:24]   = Image[374];
    assign  image_0_320[23:16]   = Image[404];
    assign  image_0_320[15:8]    = Image[405];
    assign  image_0_320[7:0]     = Image[406];

    assign  image_0_321[71:64]   = Image[341];
    assign  image_0_321[63:56]   = Image[342];
    assign  image_0_321[55:48]   = Image[343];
    assign  image_0_321[47:40]   = Image[373];
    assign  image_0_321[39:32]   = Image[374];
    assign  image_0_321[31:24]   = Image[375];
    assign  image_0_321[23:16]   = Image[405];
    assign  image_0_321[15:8]    = Image[406];
    assign  image_0_321[7:0]     = Image[407];

    assign  image_0_322[71:64]   = Image[342];
    assign  image_0_322[63:56]   = Image[343];
    assign  image_0_322[55:48]   = Image[344];
    assign  image_0_322[47:40]   = Image[374];
    assign  image_0_322[39:32]   = Image[375];
    assign  image_0_322[31:24]   = Image[376];
    assign  image_0_322[23:16]   = Image[406];
    assign  image_0_322[15:8]    = Image[407];
    assign  image_0_322[7:0]     = Image[408];

    assign  image_0_323[71:64]   = Image[343];
    assign  image_0_323[63:56]   = Image[344];
    assign  image_0_323[55:48]   = Image[345];
    assign  image_0_323[47:40]   = Image[375];
    assign  image_0_323[39:32]   = Image[376];
    assign  image_0_323[31:24]   = Image[377];
    assign  image_0_323[23:16]   = Image[407];
    assign  image_0_323[15:8]    = Image[408];
    assign  image_0_323[7:0]     = Image[409];

    assign  image_0_324[71:64]   = Image[344];
    assign  image_0_324[63:56]   = Image[345];
    assign  image_0_324[55:48]   = Image[346];
    assign  image_0_324[47:40]   = Image[376];
    assign  image_0_324[39:32]   = Image[377];
    assign  image_0_324[31:24]   = Image[378];
    assign  image_0_324[23:16]   = Image[408];
    assign  image_0_324[15:8]    = Image[409];
    assign  image_0_324[7:0]     = Image[410];

    assign  image_0_325[71:64]   = Image[345];
    assign  image_0_325[63:56]   = Image[346];
    assign  image_0_325[55:48]   = Image[347];
    assign  image_0_325[47:40]   = Image[377];
    assign  image_0_325[39:32]   = Image[378];
    assign  image_0_325[31:24]   = Image[379];
    assign  image_0_325[23:16]   = Image[409];
    assign  image_0_325[15:8]    = Image[410];
    assign  image_0_325[7:0]     = Image[411];

    assign  image_0_326[71:64]   = Image[346];
    assign  image_0_326[63:56]   = Image[347];
    assign  image_0_326[55:48]   = Image[348];
    assign  image_0_326[47:40]   = Image[378];
    assign  image_0_326[39:32]   = Image[379];
    assign  image_0_326[31:24]   = Image[380];
    assign  image_0_326[23:16]   = Image[410];
    assign  image_0_326[15:8]    = Image[411];
    assign  image_0_326[7:0]     = Image[412];

    assign  image_0_327[71:64]   = Image[347];
    assign  image_0_327[63:56]   = Image[348];
    assign  image_0_327[55:48]   = Image[349];
    assign  image_0_327[47:40]   = Image[379];
    assign  image_0_327[39:32]   = Image[380];
    assign  image_0_327[31:24]   = Image[381];
    assign  image_0_327[23:16]   = Image[411];
    assign  image_0_327[15:8]    = Image[412];
    assign  image_0_327[7:0]     = Image[413];

    assign  image_0_328[71:64]   = Image[348];
    assign  image_0_328[63:56]   = Image[349];
    assign  image_0_328[55:48]   = Image[350];
    assign  image_0_328[47:40]   = Image[380];
    assign  image_0_328[39:32]   = Image[381];
    assign  image_0_328[31:24]   = Image[382];
    assign  image_0_328[23:16]   = Image[412];
    assign  image_0_328[15:8]    = Image[413];
    assign  image_0_328[7:0]     = Image[414];

    assign  image_0_329[71:64]   = Image[349];
    assign  image_0_329[63:56]   = Image[350];
    assign  image_0_329[55:48]   = Image[351];
    assign  image_0_329[47:40]   = Image[381];
    assign  image_0_329[39:32]   = Image[382];
    assign  image_0_329[31:24]   = Image[383];
    assign  image_0_329[23:16]   = Image[413];
    assign  image_0_329[15:8]    = Image[414];
    assign  image_0_329[7:0]     = Image[415];

    assign  image_0_330[71:64]   = Image[352];
    assign  image_0_330[63:56]   = Image[353];
    assign  image_0_330[55:48]   = Image[354];
    assign  image_0_330[47:40]   = Image[384];
    assign  image_0_330[39:32]   = Image[385];
    assign  image_0_330[31:24]   = Image[386];
    assign  image_0_330[23:16]   = Image[416];
    assign  image_0_330[15:8]    = Image[417];
    assign  image_0_330[7:0]     = Image[418];

    assign  image_0_331[71:64]   = Image[353];
    assign  image_0_331[63:56]   = Image[354];
    assign  image_0_331[55:48]   = Image[355];
    assign  image_0_331[47:40]   = Image[385];
    assign  image_0_331[39:32]   = Image[386];
    assign  image_0_331[31:24]   = Image[387];
    assign  image_0_331[23:16]   = Image[417];
    assign  image_0_331[15:8]    = Image[418];
    assign  image_0_331[7:0]     = Image[419];

    assign  image_0_332[71:64]   = Image[354];
    assign  image_0_332[63:56]   = Image[355];
    assign  image_0_332[55:48]   = Image[356];
    assign  image_0_332[47:40]   = Image[386];
    assign  image_0_332[39:32]   = Image[387];
    assign  image_0_332[31:24]   = Image[388];
    assign  image_0_332[23:16]   = Image[418];
    assign  image_0_332[15:8]    = Image[419];
    assign  image_0_332[7:0]     = Image[420];

    assign  image_0_333[71:64]   = Image[355];
    assign  image_0_333[63:56]   = Image[356];
    assign  image_0_333[55:48]   = Image[357];
    assign  image_0_333[47:40]   = Image[387];
    assign  image_0_333[39:32]   = Image[388];
    assign  image_0_333[31:24]   = Image[389];
    assign  image_0_333[23:16]   = Image[419];
    assign  image_0_333[15:8]    = Image[420];
    assign  image_0_333[7:0]     = Image[421];

    assign  image_0_334[71:64]   = Image[356];
    assign  image_0_334[63:56]   = Image[357];
    assign  image_0_334[55:48]   = Image[358];
    assign  image_0_334[47:40]   = Image[388];
    assign  image_0_334[39:32]   = Image[389];
    assign  image_0_334[31:24]   = Image[390];
    assign  image_0_334[23:16]   = Image[420];
    assign  image_0_334[15:8]    = Image[421];
    assign  image_0_334[7:0]     = Image[422];

    assign  image_0_335[71:64]   = Image[357];
    assign  image_0_335[63:56]   = Image[358];
    assign  image_0_335[55:48]   = Image[359];
    assign  image_0_335[47:40]   = Image[389];
    assign  image_0_335[39:32]   = Image[390];
    assign  image_0_335[31:24]   = Image[391];
    assign  image_0_335[23:16]   = Image[421];
    assign  image_0_335[15:8]    = Image[422];
    assign  image_0_335[7:0]     = Image[423];

    assign  image_0_336[71:64]   = Image[358];
    assign  image_0_336[63:56]   = Image[359];
    assign  image_0_336[55:48]   = Image[360];
    assign  image_0_336[47:40]   = Image[390];
    assign  image_0_336[39:32]   = Image[391];
    assign  image_0_336[31:24]   = Image[392];
    assign  image_0_336[23:16]   = Image[422];
    assign  image_0_336[15:8]    = Image[423];
    assign  image_0_336[7:0]     = Image[424];

    assign  image_0_337[71:64]   = Image[359];
    assign  image_0_337[63:56]   = Image[360];
    assign  image_0_337[55:48]   = Image[361];
    assign  image_0_337[47:40]   = Image[391];
    assign  image_0_337[39:32]   = Image[392];
    assign  image_0_337[31:24]   = Image[393];
    assign  image_0_337[23:16]   = Image[423];
    assign  image_0_337[15:8]    = Image[424];
    assign  image_0_337[7:0]     = Image[425];

    assign  image_0_338[71:64]   = Image[360];
    assign  image_0_338[63:56]   = Image[361];
    assign  image_0_338[55:48]   = Image[362];
    assign  image_0_338[47:40]   = Image[392];
    assign  image_0_338[39:32]   = Image[393];
    assign  image_0_338[31:24]   = Image[394];
    assign  image_0_338[23:16]   = Image[424];
    assign  image_0_338[15:8]    = Image[425];
    assign  image_0_338[7:0]     = Image[426];

    assign  image_0_339[71:64]   = Image[361];
    assign  image_0_339[63:56]   = Image[362];
    assign  image_0_339[55:48]   = Image[363];
    assign  image_0_339[47:40]   = Image[393];
    assign  image_0_339[39:32]   = Image[394];
    assign  image_0_339[31:24]   = Image[395];
    assign  image_0_339[23:16]   = Image[425];
    assign  image_0_339[15:8]    = Image[426];
    assign  image_0_339[7:0]     = Image[427];

    assign  image_0_340[71:64]   = Image[362];
    assign  image_0_340[63:56]   = Image[363];
    assign  image_0_340[55:48]   = Image[364];
    assign  image_0_340[47:40]   = Image[394];
    assign  image_0_340[39:32]   = Image[395];
    assign  image_0_340[31:24]   = Image[396];
    assign  image_0_340[23:16]   = Image[426];
    assign  image_0_340[15:8]    = Image[427];
    assign  image_0_340[7:0]     = Image[428];

    assign  image_0_341[71:64]   = Image[363];
    assign  image_0_341[63:56]   = Image[364];
    assign  image_0_341[55:48]   = Image[365];
    assign  image_0_341[47:40]   = Image[395];
    assign  image_0_341[39:32]   = Image[396];
    assign  image_0_341[31:24]   = Image[397];
    assign  image_0_341[23:16]   = Image[427];
    assign  image_0_341[15:8]    = Image[428];
    assign  image_0_341[7:0]     = Image[429];

    assign  image_0_342[71:64]   = Image[364];
    assign  image_0_342[63:56]   = Image[365];
    assign  image_0_342[55:48]   = Image[366];
    assign  image_0_342[47:40]   = Image[396];
    assign  image_0_342[39:32]   = Image[397];
    assign  image_0_342[31:24]   = Image[398];
    assign  image_0_342[23:16]   = Image[428];
    assign  image_0_342[15:8]    = Image[429];
    assign  image_0_342[7:0]     = Image[430];

    assign  image_0_343[71:64]   = Image[365];
    assign  image_0_343[63:56]   = Image[366];
    assign  image_0_343[55:48]   = Image[367];
    assign  image_0_343[47:40]   = Image[397];
    assign  image_0_343[39:32]   = Image[398];
    assign  image_0_343[31:24]   = Image[399];
    assign  image_0_343[23:16]   = Image[429];
    assign  image_0_343[15:8]    = Image[430];
    assign  image_0_343[7:0]     = Image[431];

    assign  image_0_344[71:64]   = Image[366];
    assign  image_0_344[63:56]   = Image[367];
    assign  image_0_344[55:48]   = Image[368];
    assign  image_0_344[47:40]   = Image[398];
    assign  image_0_344[39:32]   = Image[399];
    assign  image_0_344[31:24]   = Image[400];
    assign  image_0_344[23:16]   = Image[430];
    assign  image_0_344[15:8]    = Image[431];
    assign  image_0_344[7:0]     = Image[432];

    assign  image_0_345[71:64]   = Image[367];
    assign  image_0_345[63:56]   = Image[368];
    assign  image_0_345[55:48]   = Image[369];
    assign  image_0_345[47:40]   = Image[399];
    assign  image_0_345[39:32]   = Image[400];
    assign  image_0_345[31:24]   = Image[401];
    assign  image_0_345[23:16]   = Image[431];
    assign  image_0_345[15:8]    = Image[432];
    assign  image_0_345[7:0]     = Image[433];

    assign  image_0_346[71:64]   = Image[368];
    assign  image_0_346[63:56]   = Image[369];
    assign  image_0_346[55:48]   = Image[370];
    assign  image_0_346[47:40]   = Image[400];
    assign  image_0_346[39:32]   = Image[401];
    assign  image_0_346[31:24]   = Image[402];
    assign  image_0_346[23:16]   = Image[432];
    assign  image_0_346[15:8]    = Image[433];
    assign  image_0_346[7:0]     = Image[434];

    assign  image_0_347[71:64]   = Image[369];
    assign  image_0_347[63:56]   = Image[370];
    assign  image_0_347[55:48]   = Image[371];
    assign  image_0_347[47:40]   = Image[401];
    assign  image_0_347[39:32]   = Image[402];
    assign  image_0_347[31:24]   = Image[403];
    assign  image_0_347[23:16]   = Image[433];
    assign  image_0_347[15:8]    = Image[434];
    assign  image_0_347[7:0]     = Image[435];

    assign  image_0_348[71:64]   = Image[370];
    assign  image_0_348[63:56]   = Image[371];
    assign  image_0_348[55:48]   = Image[372];
    assign  image_0_348[47:40]   = Image[402];
    assign  image_0_348[39:32]   = Image[403];
    assign  image_0_348[31:24]   = Image[404];
    assign  image_0_348[23:16]   = Image[434];
    assign  image_0_348[15:8]    = Image[435];
    assign  image_0_348[7:0]     = Image[436];

    assign  image_0_349[71:64]   = Image[371];
    assign  image_0_349[63:56]   = Image[372];
    assign  image_0_349[55:48]   = Image[373];
    assign  image_0_349[47:40]   = Image[403];
    assign  image_0_349[39:32]   = Image[404];
    assign  image_0_349[31:24]   = Image[405];
    assign  image_0_349[23:16]   = Image[435];
    assign  image_0_349[15:8]    = Image[436];
    assign  image_0_349[7:0]     = Image[437];

    assign  image_0_350[71:64]   = Image[372];
    assign  image_0_350[63:56]   = Image[373];
    assign  image_0_350[55:48]   = Image[374];
    assign  image_0_350[47:40]   = Image[404];
    assign  image_0_350[39:32]   = Image[405];
    assign  image_0_350[31:24]   = Image[406];
    assign  image_0_350[23:16]   = Image[436];
    assign  image_0_350[15:8]    = Image[437];
    assign  image_0_350[7:0]     = Image[438];

    assign  image_0_351[71:64]   = Image[373];
    assign  image_0_351[63:56]   = Image[374];
    assign  image_0_351[55:48]   = Image[375];
    assign  image_0_351[47:40]   = Image[405];
    assign  image_0_351[39:32]   = Image[406];
    assign  image_0_351[31:24]   = Image[407];
    assign  image_0_351[23:16]   = Image[437];
    assign  image_0_351[15:8]    = Image[438];
    assign  image_0_351[7:0]     = Image[439];

    assign  image_0_352[71:64]   = Image[374];
    assign  image_0_352[63:56]   = Image[375];
    assign  image_0_352[55:48]   = Image[376];
    assign  image_0_352[47:40]   = Image[406];
    assign  image_0_352[39:32]   = Image[407];
    assign  image_0_352[31:24]   = Image[408];
    assign  image_0_352[23:16]   = Image[438];
    assign  image_0_352[15:8]    = Image[439];
    assign  image_0_352[7:0]     = Image[440];

    assign  image_0_353[71:64]   = Image[375];
    assign  image_0_353[63:56]   = Image[376];
    assign  image_0_353[55:48]   = Image[377];
    assign  image_0_353[47:40]   = Image[407];
    assign  image_0_353[39:32]   = Image[408];
    assign  image_0_353[31:24]   = Image[409];
    assign  image_0_353[23:16]   = Image[439];
    assign  image_0_353[15:8]    = Image[440];
    assign  image_0_353[7:0]     = Image[441];

    assign  image_0_354[71:64]   = Image[376];
    assign  image_0_354[63:56]   = Image[377];
    assign  image_0_354[55:48]   = Image[378];
    assign  image_0_354[47:40]   = Image[408];
    assign  image_0_354[39:32]   = Image[409];
    assign  image_0_354[31:24]   = Image[410];
    assign  image_0_354[23:16]   = Image[440];
    assign  image_0_354[15:8]    = Image[441];
    assign  image_0_354[7:0]     = Image[442];

    assign  image_0_355[71:64]   = Image[377];
    assign  image_0_355[63:56]   = Image[378];
    assign  image_0_355[55:48]   = Image[379];
    assign  image_0_355[47:40]   = Image[409];
    assign  image_0_355[39:32]   = Image[410];
    assign  image_0_355[31:24]   = Image[411];
    assign  image_0_355[23:16]   = Image[441];
    assign  image_0_355[15:8]    = Image[442];
    assign  image_0_355[7:0]     = Image[443];

    assign  image_0_356[71:64]   = Image[378];
    assign  image_0_356[63:56]   = Image[379];
    assign  image_0_356[55:48]   = Image[380];
    assign  image_0_356[47:40]   = Image[410];
    assign  image_0_356[39:32]   = Image[411];
    assign  image_0_356[31:24]   = Image[412];
    assign  image_0_356[23:16]   = Image[442];
    assign  image_0_356[15:8]    = Image[443];
    assign  image_0_356[7:0]     = Image[444];

    assign  image_0_357[71:64]   = Image[379];
    assign  image_0_357[63:56]   = Image[380];
    assign  image_0_357[55:48]   = Image[381];
    assign  image_0_357[47:40]   = Image[411];
    assign  image_0_357[39:32]   = Image[412];
    assign  image_0_357[31:24]   = Image[413];
    assign  image_0_357[23:16]   = Image[443];
    assign  image_0_357[15:8]    = Image[444];
    assign  image_0_357[7:0]     = Image[445];

    assign  image_0_358[71:64]   = Image[380];
    assign  image_0_358[63:56]   = Image[381];
    assign  image_0_358[55:48]   = Image[382];
    assign  image_0_358[47:40]   = Image[412];
    assign  image_0_358[39:32]   = Image[413];
    assign  image_0_358[31:24]   = Image[414];
    assign  image_0_358[23:16]   = Image[444];
    assign  image_0_358[15:8]    = Image[445];
    assign  image_0_358[7:0]     = Image[446];

    assign  image_0_359[71:64]   = Image[381];
    assign  image_0_359[63:56]   = Image[382];
    assign  image_0_359[55:48]   = Image[383];
    assign  image_0_359[47:40]   = Image[413];
    assign  image_0_359[39:32]   = Image[414];
    assign  image_0_359[31:24]   = Image[415];
    assign  image_0_359[23:16]   = Image[445];
    assign  image_0_359[15:8]    = Image[446];
    assign  image_0_359[7:0]     = Image[447];

    assign  image_0_360[71:64]   = Image[384];
    assign  image_0_360[63:56]   = Image[385];
    assign  image_0_360[55:48]   = Image[386];
    assign  image_0_360[47:40]   = Image[416];
    assign  image_0_360[39:32]   = Image[417];
    assign  image_0_360[31:24]   = Image[418];
    assign  image_0_360[23:16]   = Image[448];
    assign  image_0_360[15:8]    = Image[449];
    assign  image_0_360[7:0]     = Image[450];

    assign  image_0_361[71:64]   = Image[385];
    assign  image_0_361[63:56]   = Image[386];
    assign  image_0_361[55:48]   = Image[387];
    assign  image_0_361[47:40]   = Image[417];
    assign  image_0_361[39:32]   = Image[418];
    assign  image_0_361[31:24]   = Image[419];
    assign  image_0_361[23:16]   = Image[449];
    assign  image_0_361[15:8]    = Image[450];
    assign  image_0_361[7:0]     = Image[451];

    assign  image_0_362[71:64]   = Image[386];
    assign  image_0_362[63:56]   = Image[387];
    assign  image_0_362[55:48]   = Image[388];
    assign  image_0_362[47:40]   = Image[418];
    assign  image_0_362[39:32]   = Image[419];
    assign  image_0_362[31:24]   = Image[420];
    assign  image_0_362[23:16]   = Image[450];
    assign  image_0_362[15:8]    = Image[451];
    assign  image_0_362[7:0]     = Image[452];

    assign  image_0_363[71:64]   = Image[387];
    assign  image_0_363[63:56]   = Image[388];
    assign  image_0_363[55:48]   = Image[389];
    assign  image_0_363[47:40]   = Image[419];
    assign  image_0_363[39:32]   = Image[420];
    assign  image_0_363[31:24]   = Image[421];
    assign  image_0_363[23:16]   = Image[451];
    assign  image_0_363[15:8]    = Image[452];
    assign  image_0_363[7:0]     = Image[453];

    assign  image_0_364[71:64]   = Image[388];
    assign  image_0_364[63:56]   = Image[389];
    assign  image_0_364[55:48]   = Image[390];
    assign  image_0_364[47:40]   = Image[420];
    assign  image_0_364[39:32]   = Image[421];
    assign  image_0_364[31:24]   = Image[422];
    assign  image_0_364[23:16]   = Image[452];
    assign  image_0_364[15:8]    = Image[453];
    assign  image_0_364[7:0]     = Image[454];

    assign  image_0_365[71:64]   = Image[389];
    assign  image_0_365[63:56]   = Image[390];
    assign  image_0_365[55:48]   = Image[391];
    assign  image_0_365[47:40]   = Image[421];
    assign  image_0_365[39:32]   = Image[422];
    assign  image_0_365[31:24]   = Image[423];
    assign  image_0_365[23:16]   = Image[453];
    assign  image_0_365[15:8]    = Image[454];
    assign  image_0_365[7:0]     = Image[455];

    assign  image_0_366[71:64]   = Image[390];
    assign  image_0_366[63:56]   = Image[391];
    assign  image_0_366[55:48]   = Image[392];
    assign  image_0_366[47:40]   = Image[422];
    assign  image_0_366[39:32]   = Image[423];
    assign  image_0_366[31:24]   = Image[424];
    assign  image_0_366[23:16]   = Image[454];
    assign  image_0_366[15:8]    = Image[455];
    assign  image_0_366[7:0]     = Image[456];

    assign  image_0_367[71:64]   = Image[391];
    assign  image_0_367[63:56]   = Image[392];
    assign  image_0_367[55:48]   = Image[393];
    assign  image_0_367[47:40]   = Image[423];
    assign  image_0_367[39:32]   = Image[424];
    assign  image_0_367[31:24]   = Image[425];
    assign  image_0_367[23:16]   = Image[455];
    assign  image_0_367[15:8]    = Image[456];
    assign  image_0_367[7:0]     = Image[457];

    assign  image_0_368[71:64]   = Image[392];
    assign  image_0_368[63:56]   = Image[393];
    assign  image_0_368[55:48]   = Image[394];
    assign  image_0_368[47:40]   = Image[424];
    assign  image_0_368[39:32]   = Image[425];
    assign  image_0_368[31:24]   = Image[426];
    assign  image_0_368[23:16]   = Image[456];
    assign  image_0_368[15:8]    = Image[457];
    assign  image_0_368[7:0]     = Image[458];

    assign  image_0_369[71:64]   = Image[393];
    assign  image_0_369[63:56]   = Image[394];
    assign  image_0_369[55:48]   = Image[395];
    assign  image_0_369[47:40]   = Image[425];
    assign  image_0_369[39:32]   = Image[426];
    assign  image_0_369[31:24]   = Image[427];
    assign  image_0_369[23:16]   = Image[457];
    assign  image_0_369[15:8]    = Image[458];
    assign  image_0_369[7:0]     = Image[459];

    assign  image_0_370[71:64]   = Image[394];
    assign  image_0_370[63:56]   = Image[395];
    assign  image_0_370[55:48]   = Image[396];
    assign  image_0_370[47:40]   = Image[426];
    assign  image_0_370[39:32]   = Image[427];
    assign  image_0_370[31:24]   = Image[428];
    assign  image_0_370[23:16]   = Image[458];
    assign  image_0_370[15:8]    = Image[459];
    assign  image_0_370[7:0]     = Image[460];

    assign  image_0_371[71:64]   = Image[395];
    assign  image_0_371[63:56]   = Image[396];
    assign  image_0_371[55:48]   = Image[397];
    assign  image_0_371[47:40]   = Image[427];
    assign  image_0_371[39:32]   = Image[428];
    assign  image_0_371[31:24]   = Image[429];
    assign  image_0_371[23:16]   = Image[459];
    assign  image_0_371[15:8]    = Image[460];
    assign  image_0_371[7:0]     = Image[461];

    assign  image_0_372[71:64]   = Image[396];
    assign  image_0_372[63:56]   = Image[397];
    assign  image_0_372[55:48]   = Image[398];
    assign  image_0_372[47:40]   = Image[428];
    assign  image_0_372[39:32]   = Image[429];
    assign  image_0_372[31:24]   = Image[430];
    assign  image_0_372[23:16]   = Image[460];
    assign  image_0_372[15:8]    = Image[461];
    assign  image_0_372[7:0]     = Image[462];

    assign  image_0_373[71:64]   = Image[397];
    assign  image_0_373[63:56]   = Image[398];
    assign  image_0_373[55:48]   = Image[399];
    assign  image_0_373[47:40]   = Image[429];
    assign  image_0_373[39:32]   = Image[430];
    assign  image_0_373[31:24]   = Image[431];
    assign  image_0_373[23:16]   = Image[461];
    assign  image_0_373[15:8]    = Image[462];
    assign  image_0_373[7:0]     = Image[463];

    assign  image_0_374[71:64]   = Image[398];
    assign  image_0_374[63:56]   = Image[399];
    assign  image_0_374[55:48]   = Image[400];
    assign  image_0_374[47:40]   = Image[430];
    assign  image_0_374[39:32]   = Image[431];
    assign  image_0_374[31:24]   = Image[432];
    assign  image_0_374[23:16]   = Image[462];
    assign  image_0_374[15:8]    = Image[463];
    assign  image_0_374[7:0]     = Image[464];

    assign  image_0_375[71:64]   = Image[399];
    assign  image_0_375[63:56]   = Image[400];
    assign  image_0_375[55:48]   = Image[401];
    assign  image_0_375[47:40]   = Image[431];
    assign  image_0_375[39:32]   = Image[432];
    assign  image_0_375[31:24]   = Image[433];
    assign  image_0_375[23:16]   = Image[463];
    assign  image_0_375[15:8]    = Image[464];
    assign  image_0_375[7:0]     = Image[465];

    assign  image_0_376[71:64]   = Image[400];
    assign  image_0_376[63:56]   = Image[401];
    assign  image_0_376[55:48]   = Image[402];
    assign  image_0_376[47:40]   = Image[432];
    assign  image_0_376[39:32]   = Image[433];
    assign  image_0_376[31:24]   = Image[434];
    assign  image_0_376[23:16]   = Image[464];
    assign  image_0_376[15:8]    = Image[465];
    assign  image_0_376[7:0]     = Image[466];

    assign  image_0_377[71:64]   = Image[401];
    assign  image_0_377[63:56]   = Image[402];
    assign  image_0_377[55:48]   = Image[403];
    assign  image_0_377[47:40]   = Image[433];
    assign  image_0_377[39:32]   = Image[434];
    assign  image_0_377[31:24]   = Image[435];
    assign  image_0_377[23:16]   = Image[465];
    assign  image_0_377[15:8]    = Image[466];
    assign  image_0_377[7:0]     = Image[467];

    assign  image_0_378[71:64]   = Image[402];
    assign  image_0_378[63:56]   = Image[403];
    assign  image_0_378[55:48]   = Image[404];
    assign  image_0_378[47:40]   = Image[434];
    assign  image_0_378[39:32]   = Image[435];
    assign  image_0_378[31:24]   = Image[436];
    assign  image_0_378[23:16]   = Image[466];
    assign  image_0_378[15:8]    = Image[467];
    assign  image_0_378[7:0]     = Image[468];

    assign  image_0_379[71:64]   = Image[403];
    assign  image_0_379[63:56]   = Image[404];
    assign  image_0_379[55:48]   = Image[405];
    assign  image_0_379[47:40]   = Image[435];
    assign  image_0_379[39:32]   = Image[436];
    assign  image_0_379[31:24]   = Image[437];
    assign  image_0_379[23:16]   = Image[467];
    assign  image_0_379[15:8]    = Image[468];
    assign  image_0_379[7:0]     = Image[469];

    assign  image_0_380[71:64]   = Image[404];
    assign  image_0_380[63:56]   = Image[405];
    assign  image_0_380[55:48]   = Image[406];
    assign  image_0_380[47:40]   = Image[436];
    assign  image_0_380[39:32]   = Image[437];
    assign  image_0_380[31:24]   = Image[438];
    assign  image_0_380[23:16]   = Image[468];
    assign  image_0_380[15:8]    = Image[469];
    assign  image_0_380[7:0]     = Image[470];

    assign  image_0_381[71:64]   = Image[405];
    assign  image_0_381[63:56]   = Image[406];
    assign  image_0_381[55:48]   = Image[407];
    assign  image_0_381[47:40]   = Image[437];
    assign  image_0_381[39:32]   = Image[438];
    assign  image_0_381[31:24]   = Image[439];
    assign  image_0_381[23:16]   = Image[469];
    assign  image_0_381[15:8]    = Image[470];
    assign  image_0_381[7:0]     = Image[471];

    assign  image_0_382[71:64]   = Image[406];
    assign  image_0_382[63:56]   = Image[407];
    assign  image_0_382[55:48]   = Image[408];
    assign  image_0_382[47:40]   = Image[438];
    assign  image_0_382[39:32]   = Image[439];
    assign  image_0_382[31:24]   = Image[440];
    assign  image_0_382[23:16]   = Image[470];
    assign  image_0_382[15:8]    = Image[471];
    assign  image_0_382[7:0]     = Image[472];

    assign  image_0_383[71:64]   = Image[407];
    assign  image_0_383[63:56]   = Image[408];
    assign  image_0_383[55:48]   = Image[409];
    assign  image_0_383[47:40]   = Image[439];
    assign  image_0_383[39:32]   = Image[440];
    assign  image_0_383[31:24]   = Image[441];
    assign  image_0_383[23:16]   = Image[471];
    assign  image_0_383[15:8]    = Image[472];
    assign  image_0_383[7:0]     = Image[473];

    assign  image_0_384[71:64]   = Image[408];
    assign  image_0_384[63:56]   = Image[409];
    assign  image_0_384[55:48]   = Image[410];
    assign  image_0_384[47:40]   = Image[440];
    assign  image_0_384[39:32]   = Image[441];
    assign  image_0_384[31:24]   = Image[442];
    assign  image_0_384[23:16]   = Image[472];
    assign  image_0_384[15:8]    = Image[473];
    assign  image_0_384[7:0]     = Image[474];

    assign  image_0_385[71:64]   = Image[409];
    assign  image_0_385[63:56]   = Image[410];
    assign  image_0_385[55:48]   = Image[411];
    assign  image_0_385[47:40]   = Image[441];
    assign  image_0_385[39:32]   = Image[442];
    assign  image_0_385[31:24]   = Image[443];
    assign  image_0_385[23:16]   = Image[473];
    assign  image_0_385[15:8]    = Image[474];
    assign  image_0_385[7:0]     = Image[475];

    assign  image_0_386[71:64]   = Image[410];
    assign  image_0_386[63:56]   = Image[411];
    assign  image_0_386[55:48]   = Image[412];
    assign  image_0_386[47:40]   = Image[442];
    assign  image_0_386[39:32]   = Image[443];
    assign  image_0_386[31:24]   = Image[444];
    assign  image_0_386[23:16]   = Image[474];
    assign  image_0_386[15:8]    = Image[475];
    assign  image_0_386[7:0]     = Image[476];

    assign  image_0_387[71:64]   = Image[411];
    assign  image_0_387[63:56]   = Image[412];
    assign  image_0_387[55:48]   = Image[413];
    assign  image_0_387[47:40]   = Image[443];
    assign  image_0_387[39:32]   = Image[444];
    assign  image_0_387[31:24]   = Image[445];
    assign  image_0_387[23:16]   = Image[475];
    assign  image_0_387[15:8]    = Image[476];
    assign  image_0_387[7:0]     = Image[477];

    assign  image_0_388[71:64]   = Image[412];
    assign  image_0_388[63:56]   = Image[413];
    assign  image_0_388[55:48]   = Image[414];
    assign  image_0_388[47:40]   = Image[444];
    assign  image_0_388[39:32]   = Image[445];
    assign  image_0_388[31:24]   = Image[446];
    assign  image_0_388[23:16]   = Image[476];
    assign  image_0_388[15:8]    = Image[477];
    assign  image_0_388[7:0]     = Image[478];

    assign  image_0_389[71:64]   = Image[413];
    assign  image_0_389[63:56]   = Image[414];
    assign  image_0_389[55:48]   = Image[415];
    assign  image_0_389[47:40]   = Image[445];
    assign  image_0_389[39:32]   = Image[446];
    assign  image_0_389[31:24]   = Image[447];
    assign  image_0_389[23:16]   = Image[477];
    assign  image_0_389[15:8]    = Image[478];
    assign  image_0_389[7:0]     = Image[479];

    assign  image_0_390[71:64]   = Image[416];
    assign  image_0_390[63:56]   = Image[417];
    assign  image_0_390[55:48]   = Image[418];
    assign  image_0_390[47:40]   = Image[448];
    assign  image_0_390[39:32]   = Image[449];
    assign  image_0_390[31:24]   = Image[450];
    assign  image_0_390[23:16]   = Image[480];
    assign  image_0_390[15:8]    = Image[481];
    assign  image_0_390[7:0]     = Image[482];

    assign  image_0_391[71:64]   = Image[417];
    assign  image_0_391[63:56]   = Image[418];
    assign  image_0_391[55:48]   = Image[419];
    assign  image_0_391[47:40]   = Image[449];
    assign  image_0_391[39:32]   = Image[450];
    assign  image_0_391[31:24]   = Image[451];
    assign  image_0_391[23:16]   = Image[481];
    assign  image_0_391[15:8]    = Image[482];
    assign  image_0_391[7:0]     = Image[483];

    assign  image_0_392[71:64]   = Image[418];
    assign  image_0_392[63:56]   = Image[419];
    assign  image_0_392[55:48]   = Image[420];
    assign  image_0_392[47:40]   = Image[450];
    assign  image_0_392[39:32]   = Image[451];
    assign  image_0_392[31:24]   = Image[452];
    assign  image_0_392[23:16]   = Image[482];
    assign  image_0_392[15:8]    = Image[483];
    assign  image_0_392[7:0]     = Image[484];

    assign  image_0_393[71:64]   = Image[419];
    assign  image_0_393[63:56]   = Image[420];
    assign  image_0_393[55:48]   = Image[421];
    assign  image_0_393[47:40]   = Image[451];
    assign  image_0_393[39:32]   = Image[452];
    assign  image_0_393[31:24]   = Image[453];
    assign  image_0_393[23:16]   = Image[483];
    assign  image_0_393[15:8]    = Image[484];
    assign  image_0_393[7:0]     = Image[485];

    assign  image_0_394[71:64]   = Image[420];
    assign  image_0_394[63:56]   = Image[421];
    assign  image_0_394[55:48]   = Image[422];
    assign  image_0_394[47:40]   = Image[452];
    assign  image_0_394[39:32]   = Image[453];
    assign  image_0_394[31:24]   = Image[454];
    assign  image_0_394[23:16]   = Image[484];
    assign  image_0_394[15:8]    = Image[485];
    assign  image_0_394[7:0]     = Image[486];

    assign  image_0_395[71:64]   = Image[421];
    assign  image_0_395[63:56]   = Image[422];
    assign  image_0_395[55:48]   = Image[423];
    assign  image_0_395[47:40]   = Image[453];
    assign  image_0_395[39:32]   = Image[454];
    assign  image_0_395[31:24]   = Image[455];
    assign  image_0_395[23:16]   = Image[485];
    assign  image_0_395[15:8]    = Image[486];
    assign  image_0_395[7:0]     = Image[487];

    assign  image_0_396[71:64]   = Image[422];
    assign  image_0_396[63:56]   = Image[423];
    assign  image_0_396[55:48]   = Image[424];
    assign  image_0_396[47:40]   = Image[454];
    assign  image_0_396[39:32]   = Image[455];
    assign  image_0_396[31:24]   = Image[456];
    assign  image_0_396[23:16]   = Image[486];
    assign  image_0_396[15:8]    = Image[487];
    assign  image_0_396[7:0]     = Image[488];

    assign  image_0_397[71:64]   = Image[423];
    assign  image_0_397[63:56]   = Image[424];
    assign  image_0_397[55:48]   = Image[425];
    assign  image_0_397[47:40]   = Image[455];
    assign  image_0_397[39:32]   = Image[456];
    assign  image_0_397[31:24]   = Image[457];
    assign  image_0_397[23:16]   = Image[487];
    assign  image_0_397[15:8]    = Image[488];
    assign  image_0_397[7:0]     = Image[489];

    assign  image_0_398[71:64]   = Image[424];
    assign  image_0_398[63:56]   = Image[425];
    assign  image_0_398[55:48]   = Image[426];
    assign  image_0_398[47:40]   = Image[456];
    assign  image_0_398[39:32]   = Image[457];
    assign  image_0_398[31:24]   = Image[458];
    assign  image_0_398[23:16]   = Image[488];
    assign  image_0_398[15:8]    = Image[489];
    assign  image_0_398[7:0]     = Image[490];

    assign  image_0_399[71:64]   = Image[425];
    assign  image_0_399[63:56]   = Image[426];
    assign  image_0_399[55:48]   = Image[427];
    assign  image_0_399[47:40]   = Image[457];
    assign  image_0_399[39:32]   = Image[458];
    assign  image_0_399[31:24]   = Image[459];
    assign  image_0_399[23:16]   = Image[489];
    assign  image_0_399[15:8]    = Image[490];
    assign  image_0_399[7:0]     = Image[491];

    assign  image_0_400[71:64]   = Image[426];
    assign  image_0_400[63:56]   = Image[427];
    assign  image_0_400[55:48]   = Image[428];
    assign  image_0_400[47:40]   = Image[458];
    assign  image_0_400[39:32]   = Image[459];
    assign  image_0_400[31:24]   = Image[460];
    assign  image_0_400[23:16]   = Image[490];
    assign  image_0_400[15:8]    = Image[491];
    assign  image_0_400[7:0]     = Image[492];

    assign  image_0_401[71:64]   = Image[427];
    assign  image_0_401[63:56]   = Image[428];
    assign  image_0_401[55:48]   = Image[429];
    assign  image_0_401[47:40]   = Image[459];
    assign  image_0_401[39:32]   = Image[460];
    assign  image_0_401[31:24]   = Image[461];
    assign  image_0_401[23:16]   = Image[491];
    assign  image_0_401[15:8]    = Image[492];
    assign  image_0_401[7:0]     = Image[493];

    assign  image_0_402[71:64]   = Image[428];
    assign  image_0_402[63:56]   = Image[429];
    assign  image_0_402[55:48]   = Image[430];
    assign  image_0_402[47:40]   = Image[460];
    assign  image_0_402[39:32]   = Image[461];
    assign  image_0_402[31:24]   = Image[462];
    assign  image_0_402[23:16]   = Image[492];
    assign  image_0_402[15:8]    = Image[493];
    assign  image_0_402[7:0]     = Image[494];

    assign  image_0_403[71:64]   = Image[429];
    assign  image_0_403[63:56]   = Image[430];
    assign  image_0_403[55:48]   = Image[431];
    assign  image_0_403[47:40]   = Image[461];
    assign  image_0_403[39:32]   = Image[462];
    assign  image_0_403[31:24]   = Image[463];
    assign  image_0_403[23:16]   = Image[493];
    assign  image_0_403[15:8]    = Image[494];
    assign  image_0_403[7:0]     = Image[495];

    assign  image_0_404[71:64]   = Image[430];
    assign  image_0_404[63:56]   = Image[431];
    assign  image_0_404[55:48]   = Image[432];
    assign  image_0_404[47:40]   = Image[462];
    assign  image_0_404[39:32]   = Image[463];
    assign  image_0_404[31:24]   = Image[464];
    assign  image_0_404[23:16]   = Image[494];
    assign  image_0_404[15:8]    = Image[495];
    assign  image_0_404[7:0]     = Image[496];

    assign  image_0_405[71:64]   = Image[431];
    assign  image_0_405[63:56]   = Image[432];
    assign  image_0_405[55:48]   = Image[433];
    assign  image_0_405[47:40]   = Image[463];
    assign  image_0_405[39:32]   = Image[464];
    assign  image_0_405[31:24]   = Image[465];
    assign  image_0_405[23:16]   = Image[495];
    assign  image_0_405[15:8]    = Image[496];
    assign  image_0_405[7:0]     = Image[497];

    assign  image_0_406[71:64]   = Image[432];
    assign  image_0_406[63:56]   = Image[433];
    assign  image_0_406[55:48]   = Image[434];
    assign  image_0_406[47:40]   = Image[464];
    assign  image_0_406[39:32]   = Image[465];
    assign  image_0_406[31:24]   = Image[466];
    assign  image_0_406[23:16]   = Image[496];
    assign  image_0_406[15:8]    = Image[497];
    assign  image_0_406[7:0]     = Image[498];

    assign  image_0_407[71:64]   = Image[433];
    assign  image_0_407[63:56]   = Image[434];
    assign  image_0_407[55:48]   = Image[435];
    assign  image_0_407[47:40]   = Image[465];
    assign  image_0_407[39:32]   = Image[466];
    assign  image_0_407[31:24]   = Image[467];
    assign  image_0_407[23:16]   = Image[497];
    assign  image_0_407[15:8]    = Image[498];
    assign  image_0_407[7:0]     = Image[499];

    assign  image_0_408[71:64]   = Image[434];
    assign  image_0_408[63:56]   = Image[435];
    assign  image_0_408[55:48]   = Image[436];
    assign  image_0_408[47:40]   = Image[466];
    assign  image_0_408[39:32]   = Image[467];
    assign  image_0_408[31:24]   = Image[468];
    assign  image_0_408[23:16]   = Image[498];
    assign  image_0_408[15:8]    = Image[499];
    assign  image_0_408[7:0]     = Image[500];

    assign  image_0_409[71:64]   = Image[435];
    assign  image_0_409[63:56]   = Image[436];
    assign  image_0_409[55:48]   = Image[437];
    assign  image_0_409[47:40]   = Image[467];
    assign  image_0_409[39:32]   = Image[468];
    assign  image_0_409[31:24]   = Image[469];
    assign  image_0_409[23:16]   = Image[499];
    assign  image_0_409[15:8]    = Image[500];
    assign  image_0_409[7:0]     = Image[501];

    assign  image_0_410[71:64]   = Image[436];
    assign  image_0_410[63:56]   = Image[437];
    assign  image_0_410[55:48]   = Image[438];
    assign  image_0_410[47:40]   = Image[468];
    assign  image_0_410[39:32]   = Image[469];
    assign  image_0_410[31:24]   = Image[470];
    assign  image_0_410[23:16]   = Image[500];
    assign  image_0_410[15:8]    = Image[501];
    assign  image_0_410[7:0]     = Image[502];

    assign  image_0_411[71:64]   = Image[437];
    assign  image_0_411[63:56]   = Image[438];
    assign  image_0_411[55:48]   = Image[439];
    assign  image_0_411[47:40]   = Image[469];
    assign  image_0_411[39:32]   = Image[470];
    assign  image_0_411[31:24]   = Image[471];
    assign  image_0_411[23:16]   = Image[501];
    assign  image_0_411[15:8]    = Image[502];
    assign  image_0_411[7:0]     = Image[503];

    assign  image_0_412[71:64]   = Image[438];
    assign  image_0_412[63:56]   = Image[439];
    assign  image_0_412[55:48]   = Image[440];
    assign  image_0_412[47:40]   = Image[470];
    assign  image_0_412[39:32]   = Image[471];
    assign  image_0_412[31:24]   = Image[472];
    assign  image_0_412[23:16]   = Image[502];
    assign  image_0_412[15:8]    = Image[503];
    assign  image_0_412[7:0]     = Image[504];

    assign  image_0_413[71:64]   = Image[439];
    assign  image_0_413[63:56]   = Image[440];
    assign  image_0_413[55:48]   = Image[441];
    assign  image_0_413[47:40]   = Image[471];
    assign  image_0_413[39:32]   = Image[472];
    assign  image_0_413[31:24]   = Image[473];
    assign  image_0_413[23:16]   = Image[503];
    assign  image_0_413[15:8]    = Image[504];
    assign  image_0_413[7:0]     = Image[505];

    assign  image_0_414[71:64]   = Image[440];
    assign  image_0_414[63:56]   = Image[441];
    assign  image_0_414[55:48]   = Image[442];
    assign  image_0_414[47:40]   = Image[472];
    assign  image_0_414[39:32]   = Image[473];
    assign  image_0_414[31:24]   = Image[474];
    assign  image_0_414[23:16]   = Image[504];
    assign  image_0_414[15:8]    = Image[505];
    assign  image_0_414[7:0]     = Image[506];

    assign  image_0_415[71:64]   = Image[441];
    assign  image_0_415[63:56]   = Image[442];
    assign  image_0_415[55:48]   = Image[443];
    assign  image_0_415[47:40]   = Image[473];
    assign  image_0_415[39:32]   = Image[474];
    assign  image_0_415[31:24]   = Image[475];
    assign  image_0_415[23:16]   = Image[505];
    assign  image_0_415[15:8]    = Image[506];
    assign  image_0_415[7:0]     = Image[507];

    assign  image_0_416[71:64]   = Image[442];
    assign  image_0_416[63:56]   = Image[443];
    assign  image_0_416[55:48]   = Image[444];
    assign  image_0_416[47:40]   = Image[474];
    assign  image_0_416[39:32]   = Image[475];
    assign  image_0_416[31:24]   = Image[476];
    assign  image_0_416[23:16]   = Image[506];
    assign  image_0_416[15:8]    = Image[507];
    assign  image_0_416[7:0]     = Image[508];

    assign  image_0_417[71:64]   = Image[443];
    assign  image_0_417[63:56]   = Image[444];
    assign  image_0_417[55:48]   = Image[445];
    assign  image_0_417[47:40]   = Image[475];
    assign  image_0_417[39:32]   = Image[476];
    assign  image_0_417[31:24]   = Image[477];
    assign  image_0_417[23:16]   = Image[507];
    assign  image_0_417[15:8]    = Image[508];
    assign  image_0_417[7:0]     = Image[509];

    assign  image_0_418[71:64]   = Image[444];
    assign  image_0_418[63:56]   = Image[445];
    assign  image_0_418[55:48]   = Image[446];
    assign  image_0_418[47:40]   = Image[476];
    assign  image_0_418[39:32]   = Image[477];
    assign  image_0_418[31:24]   = Image[478];
    assign  image_0_418[23:16]   = Image[508];
    assign  image_0_418[15:8]    = Image[509];
    assign  image_0_418[7:0]     = Image[510];

    assign  image_0_419[71:64]   = Image[445];
    assign  image_0_419[63:56]   = Image[446];
    assign  image_0_419[55:48]   = Image[447];
    assign  image_0_419[47:40]   = Image[477];
    assign  image_0_419[39:32]   = Image[478];
    assign  image_0_419[31:24]   = Image[479];
    assign  image_0_419[23:16]   = Image[509];
    assign  image_0_419[15:8]    = Image[510];
    assign  image_0_419[7:0]     = Image[511];

    assign  image_0_420[71:64]   = Image[448];
    assign  image_0_420[63:56]   = Image[449];
    assign  image_0_420[55:48]   = Image[450];
    assign  image_0_420[47:40]   = Image[480];
    assign  image_0_420[39:32]   = Image[481];
    assign  image_0_420[31:24]   = Image[482];
    assign  image_0_420[23:16]   = Image[512];
    assign  image_0_420[15:8]    = Image[513];
    assign  image_0_420[7:0]     = Image[514];

    assign  image_0_421[71:64]   = Image[449];
    assign  image_0_421[63:56]   = Image[450];
    assign  image_0_421[55:48]   = Image[451];
    assign  image_0_421[47:40]   = Image[481];
    assign  image_0_421[39:32]   = Image[482];
    assign  image_0_421[31:24]   = Image[483];
    assign  image_0_421[23:16]   = Image[513];
    assign  image_0_421[15:8]    = Image[514];
    assign  image_0_421[7:0]     = Image[515];

    assign  image_0_422[71:64]   = Image[450];
    assign  image_0_422[63:56]   = Image[451];
    assign  image_0_422[55:48]   = Image[452];
    assign  image_0_422[47:40]   = Image[482];
    assign  image_0_422[39:32]   = Image[483];
    assign  image_0_422[31:24]   = Image[484];
    assign  image_0_422[23:16]   = Image[514];
    assign  image_0_422[15:8]    = Image[515];
    assign  image_0_422[7:0]     = Image[516];

    assign  image_0_423[71:64]   = Image[451];
    assign  image_0_423[63:56]   = Image[452];
    assign  image_0_423[55:48]   = Image[453];
    assign  image_0_423[47:40]   = Image[483];
    assign  image_0_423[39:32]   = Image[484];
    assign  image_0_423[31:24]   = Image[485];
    assign  image_0_423[23:16]   = Image[515];
    assign  image_0_423[15:8]    = Image[516];
    assign  image_0_423[7:0]     = Image[517];

    assign  image_0_424[71:64]   = Image[452];
    assign  image_0_424[63:56]   = Image[453];
    assign  image_0_424[55:48]   = Image[454];
    assign  image_0_424[47:40]   = Image[484];
    assign  image_0_424[39:32]   = Image[485];
    assign  image_0_424[31:24]   = Image[486];
    assign  image_0_424[23:16]   = Image[516];
    assign  image_0_424[15:8]    = Image[517];
    assign  image_0_424[7:0]     = Image[518];

    assign  image_0_425[71:64]   = Image[453];
    assign  image_0_425[63:56]   = Image[454];
    assign  image_0_425[55:48]   = Image[455];
    assign  image_0_425[47:40]   = Image[485];
    assign  image_0_425[39:32]   = Image[486];
    assign  image_0_425[31:24]   = Image[487];
    assign  image_0_425[23:16]   = Image[517];
    assign  image_0_425[15:8]    = Image[518];
    assign  image_0_425[7:0]     = Image[519];

    assign  image_0_426[71:64]   = Image[454];
    assign  image_0_426[63:56]   = Image[455];
    assign  image_0_426[55:48]   = Image[456];
    assign  image_0_426[47:40]   = Image[486];
    assign  image_0_426[39:32]   = Image[487];
    assign  image_0_426[31:24]   = Image[488];
    assign  image_0_426[23:16]   = Image[518];
    assign  image_0_426[15:8]    = Image[519];
    assign  image_0_426[7:0]     = Image[520];

    assign  image_0_427[71:64]   = Image[455];
    assign  image_0_427[63:56]   = Image[456];
    assign  image_0_427[55:48]   = Image[457];
    assign  image_0_427[47:40]   = Image[487];
    assign  image_0_427[39:32]   = Image[488];
    assign  image_0_427[31:24]   = Image[489];
    assign  image_0_427[23:16]   = Image[519];
    assign  image_0_427[15:8]    = Image[520];
    assign  image_0_427[7:0]     = Image[521];

    assign  image_0_428[71:64]   = Image[456];
    assign  image_0_428[63:56]   = Image[457];
    assign  image_0_428[55:48]   = Image[458];
    assign  image_0_428[47:40]   = Image[488];
    assign  image_0_428[39:32]   = Image[489];
    assign  image_0_428[31:24]   = Image[490];
    assign  image_0_428[23:16]   = Image[520];
    assign  image_0_428[15:8]    = Image[521];
    assign  image_0_428[7:0]     = Image[522];

    assign  image_0_429[71:64]   = Image[457];
    assign  image_0_429[63:56]   = Image[458];
    assign  image_0_429[55:48]   = Image[459];
    assign  image_0_429[47:40]   = Image[489];
    assign  image_0_429[39:32]   = Image[490];
    assign  image_0_429[31:24]   = Image[491];
    assign  image_0_429[23:16]   = Image[521];
    assign  image_0_429[15:8]    = Image[522];
    assign  image_0_429[7:0]     = Image[523];

    assign  image_0_430[71:64]   = Image[458];
    assign  image_0_430[63:56]   = Image[459];
    assign  image_0_430[55:48]   = Image[460];
    assign  image_0_430[47:40]   = Image[490];
    assign  image_0_430[39:32]   = Image[491];
    assign  image_0_430[31:24]   = Image[492];
    assign  image_0_430[23:16]   = Image[522];
    assign  image_0_430[15:8]    = Image[523];
    assign  image_0_430[7:0]     = Image[524];

    assign  image_0_431[71:64]   = Image[459];
    assign  image_0_431[63:56]   = Image[460];
    assign  image_0_431[55:48]   = Image[461];
    assign  image_0_431[47:40]   = Image[491];
    assign  image_0_431[39:32]   = Image[492];
    assign  image_0_431[31:24]   = Image[493];
    assign  image_0_431[23:16]   = Image[523];
    assign  image_0_431[15:8]    = Image[524];
    assign  image_0_431[7:0]     = Image[525];

    assign  image_0_432[71:64]   = Image[460];
    assign  image_0_432[63:56]   = Image[461];
    assign  image_0_432[55:48]   = Image[462];
    assign  image_0_432[47:40]   = Image[492];
    assign  image_0_432[39:32]   = Image[493];
    assign  image_0_432[31:24]   = Image[494];
    assign  image_0_432[23:16]   = Image[524];
    assign  image_0_432[15:8]    = Image[525];
    assign  image_0_432[7:0]     = Image[526];

    assign  image_0_433[71:64]   = Image[461];
    assign  image_0_433[63:56]   = Image[462];
    assign  image_0_433[55:48]   = Image[463];
    assign  image_0_433[47:40]   = Image[493];
    assign  image_0_433[39:32]   = Image[494];
    assign  image_0_433[31:24]   = Image[495];
    assign  image_0_433[23:16]   = Image[525];
    assign  image_0_433[15:8]    = Image[526];
    assign  image_0_433[7:0]     = Image[527];

    assign  image_0_434[71:64]   = Image[462];
    assign  image_0_434[63:56]   = Image[463];
    assign  image_0_434[55:48]   = Image[464];
    assign  image_0_434[47:40]   = Image[494];
    assign  image_0_434[39:32]   = Image[495];
    assign  image_0_434[31:24]   = Image[496];
    assign  image_0_434[23:16]   = Image[526];
    assign  image_0_434[15:8]    = Image[527];
    assign  image_0_434[7:0]     = Image[528];

    assign  image_0_435[71:64]   = Image[463];
    assign  image_0_435[63:56]   = Image[464];
    assign  image_0_435[55:48]   = Image[465];
    assign  image_0_435[47:40]   = Image[495];
    assign  image_0_435[39:32]   = Image[496];
    assign  image_0_435[31:24]   = Image[497];
    assign  image_0_435[23:16]   = Image[527];
    assign  image_0_435[15:8]    = Image[528];
    assign  image_0_435[7:0]     = Image[529];

    assign  image_0_436[71:64]   = Image[464];
    assign  image_0_436[63:56]   = Image[465];
    assign  image_0_436[55:48]   = Image[466];
    assign  image_0_436[47:40]   = Image[496];
    assign  image_0_436[39:32]   = Image[497];
    assign  image_0_436[31:24]   = Image[498];
    assign  image_0_436[23:16]   = Image[528];
    assign  image_0_436[15:8]    = Image[529];
    assign  image_0_436[7:0]     = Image[530];

    assign  image_0_437[71:64]   = Image[465];
    assign  image_0_437[63:56]   = Image[466];
    assign  image_0_437[55:48]   = Image[467];
    assign  image_0_437[47:40]   = Image[497];
    assign  image_0_437[39:32]   = Image[498];
    assign  image_0_437[31:24]   = Image[499];
    assign  image_0_437[23:16]   = Image[529];
    assign  image_0_437[15:8]    = Image[530];
    assign  image_0_437[7:0]     = Image[531];

    assign  image_0_438[71:64]   = Image[466];
    assign  image_0_438[63:56]   = Image[467];
    assign  image_0_438[55:48]   = Image[468];
    assign  image_0_438[47:40]   = Image[498];
    assign  image_0_438[39:32]   = Image[499];
    assign  image_0_438[31:24]   = Image[500];
    assign  image_0_438[23:16]   = Image[530];
    assign  image_0_438[15:8]    = Image[531];
    assign  image_0_438[7:0]     = Image[532];

    assign  image_0_439[71:64]   = Image[467];
    assign  image_0_439[63:56]   = Image[468];
    assign  image_0_439[55:48]   = Image[469];
    assign  image_0_439[47:40]   = Image[499];
    assign  image_0_439[39:32]   = Image[500];
    assign  image_0_439[31:24]   = Image[501];
    assign  image_0_439[23:16]   = Image[531];
    assign  image_0_439[15:8]    = Image[532];
    assign  image_0_439[7:0]     = Image[533];

    assign  image_0_440[71:64]   = Image[468];
    assign  image_0_440[63:56]   = Image[469];
    assign  image_0_440[55:48]   = Image[470];
    assign  image_0_440[47:40]   = Image[500];
    assign  image_0_440[39:32]   = Image[501];
    assign  image_0_440[31:24]   = Image[502];
    assign  image_0_440[23:16]   = Image[532];
    assign  image_0_440[15:8]    = Image[533];
    assign  image_0_440[7:0]     = Image[534];

    assign  image_0_441[71:64]   = Image[469];
    assign  image_0_441[63:56]   = Image[470];
    assign  image_0_441[55:48]   = Image[471];
    assign  image_0_441[47:40]   = Image[501];
    assign  image_0_441[39:32]   = Image[502];
    assign  image_0_441[31:24]   = Image[503];
    assign  image_0_441[23:16]   = Image[533];
    assign  image_0_441[15:8]    = Image[534];
    assign  image_0_441[7:0]     = Image[535];

    assign  image_0_442[71:64]   = Image[470];
    assign  image_0_442[63:56]   = Image[471];
    assign  image_0_442[55:48]   = Image[472];
    assign  image_0_442[47:40]   = Image[502];
    assign  image_0_442[39:32]   = Image[503];
    assign  image_0_442[31:24]   = Image[504];
    assign  image_0_442[23:16]   = Image[534];
    assign  image_0_442[15:8]    = Image[535];
    assign  image_0_442[7:0]     = Image[536];

    assign  image_0_443[71:64]   = Image[471];
    assign  image_0_443[63:56]   = Image[472];
    assign  image_0_443[55:48]   = Image[473];
    assign  image_0_443[47:40]   = Image[503];
    assign  image_0_443[39:32]   = Image[504];
    assign  image_0_443[31:24]   = Image[505];
    assign  image_0_443[23:16]   = Image[535];
    assign  image_0_443[15:8]    = Image[536];
    assign  image_0_443[7:0]     = Image[537];

    assign  image_0_444[71:64]   = Image[472];
    assign  image_0_444[63:56]   = Image[473];
    assign  image_0_444[55:48]   = Image[474];
    assign  image_0_444[47:40]   = Image[504];
    assign  image_0_444[39:32]   = Image[505];
    assign  image_0_444[31:24]   = Image[506];
    assign  image_0_444[23:16]   = Image[536];
    assign  image_0_444[15:8]    = Image[537];
    assign  image_0_444[7:0]     = Image[538];

    assign  image_0_445[71:64]   = Image[473];
    assign  image_0_445[63:56]   = Image[474];
    assign  image_0_445[55:48]   = Image[475];
    assign  image_0_445[47:40]   = Image[505];
    assign  image_0_445[39:32]   = Image[506];
    assign  image_0_445[31:24]   = Image[507];
    assign  image_0_445[23:16]   = Image[537];
    assign  image_0_445[15:8]    = Image[538];
    assign  image_0_445[7:0]     = Image[539];

    assign  image_0_446[71:64]   = Image[474];
    assign  image_0_446[63:56]   = Image[475];
    assign  image_0_446[55:48]   = Image[476];
    assign  image_0_446[47:40]   = Image[506];
    assign  image_0_446[39:32]   = Image[507];
    assign  image_0_446[31:24]   = Image[508];
    assign  image_0_446[23:16]   = Image[538];
    assign  image_0_446[15:8]    = Image[539];
    assign  image_0_446[7:0]     = Image[540];

    assign  image_0_447[71:64]   = Image[475];
    assign  image_0_447[63:56]   = Image[476];
    assign  image_0_447[55:48]   = Image[477];
    assign  image_0_447[47:40]   = Image[507];
    assign  image_0_447[39:32]   = Image[508];
    assign  image_0_447[31:24]   = Image[509];
    assign  image_0_447[23:16]   = Image[539];
    assign  image_0_447[15:8]    = Image[540];
    assign  image_0_447[7:0]     = Image[541];

    assign  image_0_448[71:64]   = Image[476];
    assign  image_0_448[63:56]   = Image[477];
    assign  image_0_448[55:48]   = Image[478];
    assign  image_0_448[47:40]   = Image[508];
    assign  image_0_448[39:32]   = Image[509];
    assign  image_0_448[31:24]   = Image[510];
    assign  image_0_448[23:16]   = Image[540];
    assign  image_0_448[15:8]    = Image[541];
    assign  image_0_448[7:0]     = Image[542];

    assign  image_0_449[71:64]   = Image[477];
    assign  image_0_449[63:56]   = Image[478];
    assign  image_0_449[55:48]   = Image[479];
    assign  image_0_449[47:40]   = Image[509];
    assign  image_0_449[39:32]   = Image[510];
    assign  image_0_449[31:24]   = Image[511];
    assign  image_0_449[23:16]   = Image[541];
    assign  image_0_449[15:8]    = Image[542];
    assign  image_0_449[7:0]     = Image[543];

    assign  image_0_450[71:64]   = Image[480];
    assign  image_0_450[63:56]   = Image[481];
    assign  image_0_450[55:48]   = Image[482];
    assign  image_0_450[47:40]   = Image[512];
    assign  image_0_450[39:32]   = Image[513];
    assign  image_0_450[31:24]   = Image[514];
    assign  image_0_450[23:16]   = Image[544];
    assign  image_0_450[15:8]    = Image[545];
    assign  image_0_450[7:0]     = Image[546];

    assign  image_0_451[71:64]   = Image[481];
    assign  image_0_451[63:56]   = Image[482];
    assign  image_0_451[55:48]   = Image[483];
    assign  image_0_451[47:40]   = Image[513];
    assign  image_0_451[39:32]   = Image[514];
    assign  image_0_451[31:24]   = Image[515];
    assign  image_0_451[23:16]   = Image[545];
    assign  image_0_451[15:8]    = Image[546];
    assign  image_0_451[7:0]     = Image[547];

    assign  image_0_452[71:64]   = Image[482];
    assign  image_0_452[63:56]   = Image[483];
    assign  image_0_452[55:48]   = Image[484];
    assign  image_0_452[47:40]   = Image[514];
    assign  image_0_452[39:32]   = Image[515];
    assign  image_0_452[31:24]   = Image[516];
    assign  image_0_452[23:16]   = Image[546];
    assign  image_0_452[15:8]    = Image[547];
    assign  image_0_452[7:0]     = Image[548];

    assign  image_0_453[71:64]   = Image[483];
    assign  image_0_453[63:56]   = Image[484];
    assign  image_0_453[55:48]   = Image[485];
    assign  image_0_453[47:40]   = Image[515];
    assign  image_0_453[39:32]   = Image[516];
    assign  image_0_453[31:24]   = Image[517];
    assign  image_0_453[23:16]   = Image[547];
    assign  image_0_453[15:8]    = Image[548];
    assign  image_0_453[7:0]     = Image[549];

    assign  image_0_454[71:64]   = Image[484];
    assign  image_0_454[63:56]   = Image[485];
    assign  image_0_454[55:48]   = Image[486];
    assign  image_0_454[47:40]   = Image[516];
    assign  image_0_454[39:32]   = Image[517];
    assign  image_0_454[31:24]   = Image[518];
    assign  image_0_454[23:16]   = Image[548];
    assign  image_0_454[15:8]    = Image[549];
    assign  image_0_454[7:0]     = Image[550];

    assign  image_0_455[71:64]   = Image[485];
    assign  image_0_455[63:56]   = Image[486];
    assign  image_0_455[55:48]   = Image[487];
    assign  image_0_455[47:40]   = Image[517];
    assign  image_0_455[39:32]   = Image[518];
    assign  image_0_455[31:24]   = Image[519];
    assign  image_0_455[23:16]   = Image[549];
    assign  image_0_455[15:8]    = Image[550];
    assign  image_0_455[7:0]     = Image[551];

    assign  image_0_456[71:64]   = Image[486];
    assign  image_0_456[63:56]   = Image[487];
    assign  image_0_456[55:48]   = Image[488];
    assign  image_0_456[47:40]   = Image[518];
    assign  image_0_456[39:32]   = Image[519];
    assign  image_0_456[31:24]   = Image[520];
    assign  image_0_456[23:16]   = Image[550];
    assign  image_0_456[15:8]    = Image[551];
    assign  image_0_456[7:0]     = Image[552];

    assign  image_0_457[71:64]   = Image[487];
    assign  image_0_457[63:56]   = Image[488];
    assign  image_0_457[55:48]   = Image[489];
    assign  image_0_457[47:40]   = Image[519];
    assign  image_0_457[39:32]   = Image[520];
    assign  image_0_457[31:24]   = Image[521];
    assign  image_0_457[23:16]   = Image[551];
    assign  image_0_457[15:8]    = Image[552];
    assign  image_0_457[7:0]     = Image[553];

    assign  image_0_458[71:64]   = Image[488];
    assign  image_0_458[63:56]   = Image[489];
    assign  image_0_458[55:48]   = Image[490];
    assign  image_0_458[47:40]   = Image[520];
    assign  image_0_458[39:32]   = Image[521];
    assign  image_0_458[31:24]   = Image[522];
    assign  image_0_458[23:16]   = Image[552];
    assign  image_0_458[15:8]    = Image[553];
    assign  image_0_458[7:0]     = Image[554];

    assign  image_0_459[71:64]   = Image[489];
    assign  image_0_459[63:56]   = Image[490];
    assign  image_0_459[55:48]   = Image[491];
    assign  image_0_459[47:40]   = Image[521];
    assign  image_0_459[39:32]   = Image[522];
    assign  image_0_459[31:24]   = Image[523];
    assign  image_0_459[23:16]   = Image[553];
    assign  image_0_459[15:8]    = Image[554];
    assign  image_0_459[7:0]     = Image[555];

    assign  image_0_460[71:64]   = Image[490];
    assign  image_0_460[63:56]   = Image[491];
    assign  image_0_460[55:48]   = Image[492];
    assign  image_0_460[47:40]   = Image[522];
    assign  image_0_460[39:32]   = Image[523];
    assign  image_0_460[31:24]   = Image[524];
    assign  image_0_460[23:16]   = Image[554];
    assign  image_0_460[15:8]    = Image[555];
    assign  image_0_460[7:0]     = Image[556];

    assign  image_0_461[71:64]   = Image[491];
    assign  image_0_461[63:56]   = Image[492];
    assign  image_0_461[55:48]   = Image[493];
    assign  image_0_461[47:40]   = Image[523];
    assign  image_0_461[39:32]   = Image[524];
    assign  image_0_461[31:24]   = Image[525];
    assign  image_0_461[23:16]   = Image[555];
    assign  image_0_461[15:8]    = Image[556];
    assign  image_0_461[7:0]     = Image[557];

    assign  image_0_462[71:64]   = Image[492];
    assign  image_0_462[63:56]   = Image[493];
    assign  image_0_462[55:48]   = Image[494];
    assign  image_0_462[47:40]   = Image[524];
    assign  image_0_462[39:32]   = Image[525];
    assign  image_0_462[31:24]   = Image[526];
    assign  image_0_462[23:16]   = Image[556];
    assign  image_0_462[15:8]    = Image[557];
    assign  image_0_462[7:0]     = Image[558];

    assign  image_0_463[71:64]   = Image[493];
    assign  image_0_463[63:56]   = Image[494];
    assign  image_0_463[55:48]   = Image[495];
    assign  image_0_463[47:40]   = Image[525];
    assign  image_0_463[39:32]   = Image[526];
    assign  image_0_463[31:24]   = Image[527];
    assign  image_0_463[23:16]   = Image[557];
    assign  image_0_463[15:8]    = Image[558];
    assign  image_0_463[7:0]     = Image[559];

    assign  image_0_464[71:64]   = Image[494];
    assign  image_0_464[63:56]   = Image[495];
    assign  image_0_464[55:48]   = Image[496];
    assign  image_0_464[47:40]   = Image[526];
    assign  image_0_464[39:32]   = Image[527];
    assign  image_0_464[31:24]   = Image[528];
    assign  image_0_464[23:16]   = Image[558];
    assign  image_0_464[15:8]    = Image[559];
    assign  image_0_464[7:0]     = Image[560];

    assign  image_0_465[71:64]   = Image[495];
    assign  image_0_465[63:56]   = Image[496];
    assign  image_0_465[55:48]   = Image[497];
    assign  image_0_465[47:40]   = Image[527];
    assign  image_0_465[39:32]   = Image[528];
    assign  image_0_465[31:24]   = Image[529];
    assign  image_0_465[23:16]   = Image[559];
    assign  image_0_465[15:8]    = Image[560];
    assign  image_0_465[7:0]     = Image[561];

    assign  image_0_466[71:64]   = Image[496];
    assign  image_0_466[63:56]   = Image[497];
    assign  image_0_466[55:48]   = Image[498];
    assign  image_0_466[47:40]   = Image[528];
    assign  image_0_466[39:32]   = Image[529];
    assign  image_0_466[31:24]   = Image[530];
    assign  image_0_466[23:16]   = Image[560];
    assign  image_0_466[15:8]    = Image[561];
    assign  image_0_466[7:0]     = Image[562];

    assign  image_0_467[71:64]   = Image[497];
    assign  image_0_467[63:56]   = Image[498];
    assign  image_0_467[55:48]   = Image[499];
    assign  image_0_467[47:40]   = Image[529];
    assign  image_0_467[39:32]   = Image[530];
    assign  image_0_467[31:24]   = Image[531];
    assign  image_0_467[23:16]   = Image[561];
    assign  image_0_467[15:8]    = Image[562];
    assign  image_0_467[7:0]     = Image[563];

    assign  image_0_468[71:64]   = Image[498];
    assign  image_0_468[63:56]   = Image[499];
    assign  image_0_468[55:48]   = Image[500];
    assign  image_0_468[47:40]   = Image[530];
    assign  image_0_468[39:32]   = Image[531];
    assign  image_0_468[31:24]   = Image[532];
    assign  image_0_468[23:16]   = Image[562];
    assign  image_0_468[15:8]    = Image[563];
    assign  image_0_468[7:0]     = Image[564];

    assign  image_0_469[71:64]   = Image[499];
    assign  image_0_469[63:56]   = Image[500];
    assign  image_0_469[55:48]   = Image[501];
    assign  image_0_469[47:40]   = Image[531];
    assign  image_0_469[39:32]   = Image[532];
    assign  image_0_469[31:24]   = Image[533];
    assign  image_0_469[23:16]   = Image[563];
    assign  image_0_469[15:8]    = Image[564];
    assign  image_0_469[7:0]     = Image[565];

    assign  image_0_470[71:64]   = Image[500];
    assign  image_0_470[63:56]   = Image[501];
    assign  image_0_470[55:48]   = Image[502];
    assign  image_0_470[47:40]   = Image[532];
    assign  image_0_470[39:32]   = Image[533];
    assign  image_0_470[31:24]   = Image[534];
    assign  image_0_470[23:16]   = Image[564];
    assign  image_0_470[15:8]    = Image[565];
    assign  image_0_470[7:0]     = Image[566];

    assign  image_0_471[71:64]   = Image[501];
    assign  image_0_471[63:56]   = Image[502];
    assign  image_0_471[55:48]   = Image[503];
    assign  image_0_471[47:40]   = Image[533];
    assign  image_0_471[39:32]   = Image[534];
    assign  image_0_471[31:24]   = Image[535];
    assign  image_0_471[23:16]   = Image[565];
    assign  image_0_471[15:8]    = Image[566];
    assign  image_0_471[7:0]     = Image[567];

    assign  image_0_472[71:64]   = Image[502];
    assign  image_0_472[63:56]   = Image[503];
    assign  image_0_472[55:48]   = Image[504];
    assign  image_0_472[47:40]   = Image[534];
    assign  image_0_472[39:32]   = Image[535];
    assign  image_0_472[31:24]   = Image[536];
    assign  image_0_472[23:16]   = Image[566];
    assign  image_0_472[15:8]    = Image[567];
    assign  image_0_472[7:0]     = Image[568];

    assign  image_0_473[71:64]   = Image[503];
    assign  image_0_473[63:56]   = Image[504];
    assign  image_0_473[55:48]   = Image[505];
    assign  image_0_473[47:40]   = Image[535];
    assign  image_0_473[39:32]   = Image[536];
    assign  image_0_473[31:24]   = Image[537];
    assign  image_0_473[23:16]   = Image[567];
    assign  image_0_473[15:8]    = Image[568];
    assign  image_0_473[7:0]     = Image[569];

    assign  image_0_474[71:64]   = Image[504];
    assign  image_0_474[63:56]   = Image[505];
    assign  image_0_474[55:48]   = Image[506];
    assign  image_0_474[47:40]   = Image[536];
    assign  image_0_474[39:32]   = Image[537];
    assign  image_0_474[31:24]   = Image[538];
    assign  image_0_474[23:16]   = Image[568];
    assign  image_0_474[15:8]    = Image[569];
    assign  image_0_474[7:0]     = Image[570];

    assign  image_0_475[71:64]   = Image[505];
    assign  image_0_475[63:56]   = Image[506];
    assign  image_0_475[55:48]   = Image[507];
    assign  image_0_475[47:40]   = Image[537];
    assign  image_0_475[39:32]   = Image[538];
    assign  image_0_475[31:24]   = Image[539];
    assign  image_0_475[23:16]   = Image[569];
    assign  image_0_475[15:8]    = Image[570];
    assign  image_0_475[7:0]     = Image[571];

    assign  image_0_476[71:64]   = Image[506];
    assign  image_0_476[63:56]   = Image[507];
    assign  image_0_476[55:48]   = Image[508];
    assign  image_0_476[47:40]   = Image[538];
    assign  image_0_476[39:32]   = Image[539];
    assign  image_0_476[31:24]   = Image[540];
    assign  image_0_476[23:16]   = Image[570];
    assign  image_0_476[15:8]    = Image[571];
    assign  image_0_476[7:0]     = Image[572];

    assign  image_0_477[71:64]   = Image[507];
    assign  image_0_477[63:56]   = Image[508];
    assign  image_0_477[55:48]   = Image[509];
    assign  image_0_477[47:40]   = Image[539];
    assign  image_0_477[39:32]   = Image[540];
    assign  image_0_477[31:24]   = Image[541];
    assign  image_0_477[23:16]   = Image[571];
    assign  image_0_477[15:8]    = Image[572];
    assign  image_0_477[7:0]     = Image[573];

    assign  image_0_478[71:64]   = Image[508];
    assign  image_0_478[63:56]   = Image[509];
    assign  image_0_478[55:48]   = Image[510];
    assign  image_0_478[47:40]   = Image[540];
    assign  image_0_478[39:32]   = Image[541];
    assign  image_0_478[31:24]   = Image[542];
    assign  image_0_478[23:16]   = Image[572];
    assign  image_0_478[15:8]    = Image[573];
    assign  image_0_478[7:0]     = Image[574];

    assign  image_0_479[71:64]   = Image[509];
    assign  image_0_479[63:56]   = Image[510];
    assign  image_0_479[55:48]   = Image[511];
    assign  image_0_479[47:40]   = Image[541];
    assign  image_0_479[39:32]   = Image[542];
    assign  image_0_479[31:24]   = Image[543];
    assign  image_0_479[23:16]   = Image[573];
    assign  image_0_479[15:8]    = Image[574];
    assign  image_0_479[7:0]     = Image[575];

    assign  image_0_480[71:64]   = Image[512];
    assign  image_0_480[63:56]   = Image[513];
    assign  image_0_480[55:48]   = Image[514];
    assign  image_0_480[47:40]   = Image[544];
    assign  image_0_480[39:32]   = Image[545];
    assign  image_0_480[31:24]   = Image[546];
    assign  image_0_480[23:16]   = Image[576];
    assign  image_0_480[15:8]    = Image[577];
    assign  image_0_480[7:0]     = Image[578];

    assign  image_0_481[71:64]   = Image[513];
    assign  image_0_481[63:56]   = Image[514];
    assign  image_0_481[55:48]   = Image[515];
    assign  image_0_481[47:40]   = Image[545];
    assign  image_0_481[39:32]   = Image[546];
    assign  image_0_481[31:24]   = Image[547];
    assign  image_0_481[23:16]   = Image[577];
    assign  image_0_481[15:8]    = Image[578];
    assign  image_0_481[7:0]     = Image[579];

    assign  image_0_482[71:64]   = Image[514];
    assign  image_0_482[63:56]   = Image[515];
    assign  image_0_482[55:48]   = Image[516];
    assign  image_0_482[47:40]   = Image[546];
    assign  image_0_482[39:32]   = Image[547];
    assign  image_0_482[31:24]   = Image[548];
    assign  image_0_482[23:16]   = Image[578];
    assign  image_0_482[15:8]    = Image[579];
    assign  image_0_482[7:0]     = Image[580];

    assign  image_0_483[71:64]   = Image[515];
    assign  image_0_483[63:56]   = Image[516];
    assign  image_0_483[55:48]   = Image[517];
    assign  image_0_483[47:40]   = Image[547];
    assign  image_0_483[39:32]   = Image[548];
    assign  image_0_483[31:24]   = Image[549];
    assign  image_0_483[23:16]   = Image[579];
    assign  image_0_483[15:8]    = Image[580];
    assign  image_0_483[7:0]     = Image[581];

    assign  image_0_484[71:64]   = Image[516];
    assign  image_0_484[63:56]   = Image[517];
    assign  image_0_484[55:48]   = Image[518];
    assign  image_0_484[47:40]   = Image[548];
    assign  image_0_484[39:32]   = Image[549];
    assign  image_0_484[31:24]   = Image[550];
    assign  image_0_484[23:16]   = Image[580];
    assign  image_0_484[15:8]    = Image[581];
    assign  image_0_484[7:0]     = Image[582];

    assign  image_0_485[71:64]   = Image[517];
    assign  image_0_485[63:56]   = Image[518];
    assign  image_0_485[55:48]   = Image[519];
    assign  image_0_485[47:40]   = Image[549];
    assign  image_0_485[39:32]   = Image[550];
    assign  image_0_485[31:24]   = Image[551];
    assign  image_0_485[23:16]   = Image[581];
    assign  image_0_485[15:8]    = Image[582];
    assign  image_0_485[7:0]     = Image[583];

    assign  image_0_486[71:64]   = Image[518];
    assign  image_0_486[63:56]   = Image[519];
    assign  image_0_486[55:48]   = Image[520];
    assign  image_0_486[47:40]   = Image[550];
    assign  image_0_486[39:32]   = Image[551];
    assign  image_0_486[31:24]   = Image[552];
    assign  image_0_486[23:16]   = Image[582];
    assign  image_0_486[15:8]    = Image[583];
    assign  image_0_486[7:0]     = Image[584];

    assign  image_0_487[71:64]   = Image[519];
    assign  image_0_487[63:56]   = Image[520];
    assign  image_0_487[55:48]   = Image[521];
    assign  image_0_487[47:40]   = Image[551];
    assign  image_0_487[39:32]   = Image[552];
    assign  image_0_487[31:24]   = Image[553];
    assign  image_0_487[23:16]   = Image[583];
    assign  image_0_487[15:8]    = Image[584];
    assign  image_0_487[7:0]     = Image[585];

    assign  image_0_488[71:64]   = Image[520];
    assign  image_0_488[63:56]   = Image[521];
    assign  image_0_488[55:48]   = Image[522];
    assign  image_0_488[47:40]   = Image[552];
    assign  image_0_488[39:32]   = Image[553];
    assign  image_0_488[31:24]   = Image[554];
    assign  image_0_488[23:16]   = Image[584];
    assign  image_0_488[15:8]    = Image[585];
    assign  image_0_488[7:0]     = Image[586];

    assign  image_0_489[71:64]   = Image[521];
    assign  image_0_489[63:56]   = Image[522];
    assign  image_0_489[55:48]   = Image[523];
    assign  image_0_489[47:40]   = Image[553];
    assign  image_0_489[39:32]   = Image[554];
    assign  image_0_489[31:24]   = Image[555];
    assign  image_0_489[23:16]   = Image[585];
    assign  image_0_489[15:8]    = Image[586];
    assign  image_0_489[7:0]     = Image[587];

    assign  image_0_490[71:64]   = Image[522];
    assign  image_0_490[63:56]   = Image[523];
    assign  image_0_490[55:48]   = Image[524];
    assign  image_0_490[47:40]   = Image[554];
    assign  image_0_490[39:32]   = Image[555];
    assign  image_0_490[31:24]   = Image[556];
    assign  image_0_490[23:16]   = Image[586];
    assign  image_0_490[15:8]    = Image[587];
    assign  image_0_490[7:0]     = Image[588];

    assign  image_0_491[71:64]   = Image[523];
    assign  image_0_491[63:56]   = Image[524];
    assign  image_0_491[55:48]   = Image[525];
    assign  image_0_491[47:40]   = Image[555];
    assign  image_0_491[39:32]   = Image[556];
    assign  image_0_491[31:24]   = Image[557];
    assign  image_0_491[23:16]   = Image[587];
    assign  image_0_491[15:8]    = Image[588];
    assign  image_0_491[7:0]     = Image[589];

    assign  image_0_492[71:64]   = Image[524];
    assign  image_0_492[63:56]   = Image[525];
    assign  image_0_492[55:48]   = Image[526];
    assign  image_0_492[47:40]   = Image[556];
    assign  image_0_492[39:32]   = Image[557];
    assign  image_0_492[31:24]   = Image[558];
    assign  image_0_492[23:16]   = Image[588];
    assign  image_0_492[15:8]    = Image[589];
    assign  image_0_492[7:0]     = Image[590];

    assign  image_0_493[71:64]   = Image[525];
    assign  image_0_493[63:56]   = Image[526];
    assign  image_0_493[55:48]   = Image[527];
    assign  image_0_493[47:40]   = Image[557];
    assign  image_0_493[39:32]   = Image[558];
    assign  image_0_493[31:24]   = Image[559];
    assign  image_0_493[23:16]   = Image[589];
    assign  image_0_493[15:8]    = Image[590];
    assign  image_0_493[7:0]     = Image[591];

    assign  image_0_494[71:64]   = Image[526];
    assign  image_0_494[63:56]   = Image[527];
    assign  image_0_494[55:48]   = Image[528];
    assign  image_0_494[47:40]   = Image[558];
    assign  image_0_494[39:32]   = Image[559];
    assign  image_0_494[31:24]   = Image[560];
    assign  image_0_494[23:16]   = Image[590];
    assign  image_0_494[15:8]    = Image[591];
    assign  image_0_494[7:0]     = Image[592];

    assign  image_0_495[71:64]   = Image[527];
    assign  image_0_495[63:56]   = Image[528];
    assign  image_0_495[55:48]   = Image[529];
    assign  image_0_495[47:40]   = Image[559];
    assign  image_0_495[39:32]   = Image[560];
    assign  image_0_495[31:24]   = Image[561];
    assign  image_0_495[23:16]   = Image[591];
    assign  image_0_495[15:8]    = Image[592];
    assign  image_0_495[7:0]     = Image[593];

    assign  image_0_496[71:64]   = Image[528];
    assign  image_0_496[63:56]   = Image[529];
    assign  image_0_496[55:48]   = Image[530];
    assign  image_0_496[47:40]   = Image[560];
    assign  image_0_496[39:32]   = Image[561];
    assign  image_0_496[31:24]   = Image[562];
    assign  image_0_496[23:16]   = Image[592];
    assign  image_0_496[15:8]    = Image[593];
    assign  image_0_496[7:0]     = Image[594];

    assign  image_0_497[71:64]   = Image[529];
    assign  image_0_497[63:56]   = Image[530];
    assign  image_0_497[55:48]   = Image[531];
    assign  image_0_497[47:40]   = Image[561];
    assign  image_0_497[39:32]   = Image[562];
    assign  image_0_497[31:24]   = Image[563];
    assign  image_0_497[23:16]   = Image[593];
    assign  image_0_497[15:8]    = Image[594];
    assign  image_0_497[7:0]     = Image[595];

    assign  image_0_498[71:64]   = Image[530];
    assign  image_0_498[63:56]   = Image[531];
    assign  image_0_498[55:48]   = Image[532];
    assign  image_0_498[47:40]   = Image[562];
    assign  image_0_498[39:32]   = Image[563];
    assign  image_0_498[31:24]   = Image[564];
    assign  image_0_498[23:16]   = Image[594];
    assign  image_0_498[15:8]    = Image[595];
    assign  image_0_498[7:0]     = Image[596];

    assign  image_0_499[71:64]   = Image[531];
    assign  image_0_499[63:56]   = Image[532];
    assign  image_0_499[55:48]   = Image[533];
    assign  image_0_499[47:40]   = Image[563];
    assign  image_0_499[39:32]   = Image[564];
    assign  image_0_499[31:24]   = Image[565];
    assign  image_0_499[23:16]   = Image[595];
    assign  image_0_499[15:8]    = Image[596];
    assign  image_0_499[7:0]     = Image[597];

    assign  image_0_500[71:64]   = Image[532];
    assign  image_0_500[63:56]   = Image[533];
    assign  image_0_500[55:48]   = Image[534];
    assign  image_0_500[47:40]   = Image[564];
    assign  image_0_500[39:32]   = Image[565];
    assign  image_0_500[31:24]   = Image[566];
    assign  image_0_500[23:16]   = Image[596];
    assign  image_0_500[15:8]    = Image[597];
    assign  image_0_500[7:0]     = Image[598];

    assign  image_0_501[71:64]   = Image[533];
    assign  image_0_501[63:56]   = Image[534];
    assign  image_0_501[55:48]   = Image[535];
    assign  image_0_501[47:40]   = Image[565];
    assign  image_0_501[39:32]   = Image[566];
    assign  image_0_501[31:24]   = Image[567];
    assign  image_0_501[23:16]   = Image[597];
    assign  image_0_501[15:8]    = Image[598];
    assign  image_0_501[7:0]     = Image[599];

    assign  image_0_502[71:64]   = Image[534];
    assign  image_0_502[63:56]   = Image[535];
    assign  image_0_502[55:48]   = Image[536];
    assign  image_0_502[47:40]   = Image[566];
    assign  image_0_502[39:32]   = Image[567];
    assign  image_0_502[31:24]   = Image[568];
    assign  image_0_502[23:16]   = Image[598];
    assign  image_0_502[15:8]    = Image[599];
    assign  image_0_502[7:0]     = Image[600];

    assign  image_0_503[71:64]   = Image[535];
    assign  image_0_503[63:56]   = Image[536];
    assign  image_0_503[55:48]   = Image[537];
    assign  image_0_503[47:40]   = Image[567];
    assign  image_0_503[39:32]   = Image[568];
    assign  image_0_503[31:24]   = Image[569];
    assign  image_0_503[23:16]   = Image[599];
    assign  image_0_503[15:8]    = Image[600];
    assign  image_0_503[7:0]     = Image[601];

    assign  image_0_504[71:64]   = Image[536];
    assign  image_0_504[63:56]   = Image[537];
    assign  image_0_504[55:48]   = Image[538];
    assign  image_0_504[47:40]   = Image[568];
    assign  image_0_504[39:32]   = Image[569];
    assign  image_0_504[31:24]   = Image[570];
    assign  image_0_504[23:16]   = Image[600];
    assign  image_0_504[15:8]    = Image[601];
    assign  image_0_504[7:0]     = Image[602];

    assign  image_0_505[71:64]   = Image[537];
    assign  image_0_505[63:56]   = Image[538];
    assign  image_0_505[55:48]   = Image[539];
    assign  image_0_505[47:40]   = Image[569];
    assign  image_0_505[39:32]   = Image[570];
    assign  image_0_505[31:24]   = Image[571];
    assign  image_0_505[23:16]   = Image[601];
    assign  image_0_505[15:8]    = Image[602];
    assign  image_0_505[7:0]     = Image[603];

    assign  image_0_506[71:64]   = Image[538];
    assign  image_0_506[63:56]   = Image[539];
    assign  image_0_506[55:48]   = Image[540];
    assign  image_0_506[47:40]   = Image[570];
    assign  image_0_506[39:32]   = Image[571];
    assign  image_0_506[31:24]   = Image[572];
    assign  image_0_506[23:16]   = Image[602];
    assign  image_0_506[15:8]    = Image[603];
    assign  image_0_506[7:0]     = Image[604];

    assign  image_0_507[71:64]   = Image[539];
    assign  image_0_507[63:56]   = Image[540];
    assign  image_0_507[55:48]   = Image[541];
    assign  image_0_507[47:40]   = Image[571];
    assign  image_0_507[39:32]   = Image[572];
    assign  image_0_507[31:24]   = Image[573];
    assign  image_0_507[23:16]   = Image[603];
    assign  image_0_507[15:8]    = Image[604];
    assign  image_0_507[7:0]     = Image[605];

    assign  image_0_508[71:64]   = Image[540];
    assign  image_0_508[63:56]   = Image[541];
    assign  image_0_508[55:48]   = Image[542];
    assign  image_0_508[47:40]   = Image[572];
    assign  image_0_508[39:32]   = Image[573];
    assign  image_0_508[31:24]   = Image[574];
    assign  image_0_508[23:16]   = Image[604];
    assign  image_0_508[15:8]    = Image[605];
    assign  image_0_508[7:0]     = Image[606];

    assign  image_0_509[71:64]   = Image[541];
    assign  image_0_509[63:56]   = Image[542];
    assign  image_0_509[55:48]   = Image[543];
    assign  image_0_509[47:40]   = Image[573];
    assign  image_0_509[39:32]   = Image[574];
    assign  image_0_509[31:24]   = Image[575];
    assign  image_0_509[23:16]   = Image[605];
    assign  image_0_509[15:8]    = Image[606];
    assign  image_0_509[7:0]     = Image[607];

    assign  image_0_510[71:64]   = Image[544];
    assign  image_0_510[63:56]   = Image[545];
    assign  image_0_510[55:48]   = Image[546];
    assign  image_0_510[47:40]   = Image[576];
    assign  image_0_510[39:32]   = Image[577];
    assign  image_0_510[31:24]   = Image[578];
    assign  image_0_510[23:16]   = Image[608];
    assign  image_0_510[15:8]    = Image[609];
    assign  image_0_510[7:0]     = Image[610];

    assign  image_0_511[71:64]   = Image[545];
    assign  image_0_511[63:56]   = Image[546];
    assign  image_0_511[55:48]   = Image[547];
    assign  image_0_511[47:40]   = Image[577];
    assign  image_0_511[39:32]   = Image[578];
    assign  image_0_511[31:24]   = Image[579];
    assign  image_0_511[23:16]   = Image[609];
    assign  image_0_511[15:8]    = Image[610];
    assign  image_0_511[7:0]     = Image[611];

    assign  image_0_512[71:64]   = Image[546];
    assign  image_0_512[63:56]   = Image[547];
    assign  image_0_512[55:48]   = Image[548];
    assign  image_0_512[47:40]   = Image[578];
    assign  image_0_512[39:32]   = Image[579];
    assign  image_0_512[31:24]   = Image[580];
    assign  image_0_512[23:16]   = Image[610];
    assign  image_0_512[15:8]    = Image[611];
    assign  image_0_512[7:0]     = Image[612];

    assign  image_0_513[71:64]   = Image[547];
    assign  image_0_513[63:56]   = Image[548];
    assign  image_0_513[55:48]   = Image[549];
    assign  image_0_513[47:40]   = Image[579];
    assign  image_0_513[39:32]   = Image[580];
    assign  image_0_513[31:24]   = Image[581];
    assign  image_0_513[23:16]   = Image[611];
    assign  image_0_513[15:8]    = Image[612];
    assign  image_0_513[7:0]     = Image[613];

    assign  image_0_514[71:64]   = Image[548];
    assign  image_0_514[63:56]   = Image[549];
    assign  image_0_514[55:48]   = Image[550];
    assign  image_0_514[47:40]   = Image[580];
    assign  image_0_514[39:32]   = Image[581];
    assign  image_0_514[31:24]   = Image[582];
    assign  image_0_514[23:16]   = Image[612];
    assign  image_0_514[15:8]    = Image[613];
    assign  image_0_514[7:0]     = Image[614];

    assign  image_0_515[71:64]   = Image[549];
    assign  image_0_515[63:56]   = Image[550];
    assign  image_0_515[55:48]   = Image[551];
    assign  image_0_515[47:40]   = Image[581];
    assign  image_0_515[39:32]   = Image[582];
    assign  image_0_515[31:24]   = Image[583];
    assign  image_0_515[23:16]   = Image[613];
    assign  image_0_515[15:8]    = Image[614];
    assign  image_0_515[7:0]     = Image[615];

    assign  image_0_516[71:64]   = Image[550];
    assign  image_0_516[63:56]   = Image[551];
    assign  image_0_516[55:48]   = Image[552];
    assign  image_0_516[47:40]   = Image[582];
    assign  image_0_516[39:32]   = Image[583];
    assign  image_0_516[31:24]   = Image[584];
    assign  image_0_516[23:16]   = Image[614];
    assign  image_0_516[15:8]    = Image[615];
    assign  image_0_516[7:0]     = Image[616];

    assign  image_0_517[71:64]   = Image[551];
    assign  image_0_517[63:56]   = Image[552];
    assign  image_0_517[55:48]   = Image[553];
    assign  image_0_517[47:40]   = Image[583];
    assign  image_0_517[39:32]   = Image[584];
    assign  image_0_517[31:24]   = Image[585];
    assign  image_0_517[23:16]   = Image[615];
    assign  image_0_517[15:8]    = Image[616];
    assign  image_0_517[7:0]     = Image[617];

    assign  image_0_518[71:64]   = Image[552];
    assign  image_0_518[63:56]   = Image[553];
    assign  image_0_518[55:48]   = Image[554];
    assign  image_0_518[47:40]   = Image[584];
    assign  image_0_518[39:32]   = Image[585];
    assign  image_0_518[31:24]   = Image[586];
    assign  image_0_518[23:16]   = Image[616];
    assign  image_0_518[15:8]    = Image[617];
    assign  image_0_518[7:0]     = Image[618];

    assign  image_0_519[71:64]   = Image[553];
    assign  image_0_519[63:56]   = Image[554];
    assign  image_0_519[55:48]   = Image[555];
    assign  image_0_519[47:40]   = Image[585];
    assign  image_0_519[39:32]   = Image[586];
    assign  image_0_519[31:24]   = Image[587];
    assign  image_0_519[23:16]   = Image[617];
    assign  image_0_519[15:8]    = Image[618];
    assign  image_0_519[7:0]     = Image[619];

    assign  image_0_520[71:64]   = Image[554];
    assign  image_0_520[63:56]   = Image[555];
    assign  image_0_520[55:48]   = Image[556];
    assign  image_0_520[47:40]   = Image[586];
    assign  image_0_520[39:32]   = Image[587];
    assign  image_0_520[31:24]   = Image[588];
    assign  image_0_520[23:16]   = Image[618];
    assign  image_0_520[15:8]    = Image[619];
    assign  image_0_520[7:0]     = Image[620];

    assign  image_0_521[71:64]   = Image[555];
    assign  image_0_521[63:56]   = Image[556];
    assign  image_0_521[55:48]   = Image[557];
    assign  image_0_521[47:40]   = Image[587];
    assign  image_0_521[39:32]   = Image[588];
    assign  image_0_521[31:24]   = Image[589];
    assign  image_0_521[23:16]   = Image[619];
    assign  image_0_521[15:8]    = Image[620];
    assign  image_0_521[7:0]     = Image[621];

    assign  image_0_522[71:64]   = Image[556];
    assign  image_0_522[63:56]   = Image[557];
    assign  image_0_522[55:48]   = Image[558];
    assign  image_0_522[47:40]   = Image[588];
    assign  image_0_522[39:32]   = Image[589];
    assign  image_0_522[31:24]   = Image[590];
    assign  image_0_522[23:16]   = Image[620];
    assign  image_0_522[15:8]    = Image[621];
    assign  image_0_522[7:0]     = Image[622];

    assign  image_0_523[71:64]   = Image[557];
    assign  image_0_523[63:56]   = Image[558];
    assign  image_0_523[55:48]   = Image[559];
    assign  image_0_523[47:40]   = Image[589];
    assign  image_0_523[39:32]   = Image[590];
    assign  image_0_523[31:24]   = Image[591];
    assign  image_0_523[23:16]   = Image[621];
    assign  image_0_523[15:8]    = Image[622];
    assign  image_0_523[7:0]     = Image[623];

    assign  image_0_524[71:64]   = Image[558];
    assign  image_0_524[63:56]   = Image[559];
    assign  image_0_524[55:48]   = Image[560];
    assign  image_0_524[47:40]   = Image[590];
    assign  image_0_524[39:32]   = Image[591];
    assign  image_0_524[31:24]   = Image[592];
    assign  image_0_524[23:16]   = Image[622];
    assign  image_0_524[15:8]    = Image[623];
    assign  image_0_524[7:0]     = Image[624];

    assign  image_0_525[71:64]   = Image[559];
    assign  image_0_525[63:56]   = Image[560];
    assign  image_0_525[55:48]   = Image[561];
    assign  image_0_525[47:40]   = Image[591];
    assign  image_0_525[39:32]   = Image[592];
    assign  image_0_525[31:24]   = Image[593];
    assign  image_0_525[23:16]   = Image[623];
    assign  image_0_525[15:8]    = Image[624];
    assign  image_0_525[7:0]     = Image[625];

    assign  image_0_526[71:64]   = Image[560];
    assign  image_0_526[63:56]   = Image[561];
    assign  image_0_526[55:48]   = Image[562];
    assign  image_0_526[47:40]   = Image[592];
    assign  image_0_526[39:32]   = Image[593];
    assign  image_0_526[31:24]   = Image[594];
    assign  image_0_526[23:16]   = Image[624];
    assign  image_0_526[15:8]    = Image[625];
    assign  image_0_526[7:0]     = Image[626];

    assign  image_0_527[71:64]   = Image[561];
    assign  image_0_527[63:56]   = Image[562];
    assign  image_0_527[55:48]   = Image[563];
    assign  image_0_527[47:40]   = Image[593];
    assign  image_0_527[39:32]   = Image[594];
    assign  image_0_527[31:24]   = Image[595];
    assign  image_0_527[23:16]   = Image[625];
    assign  image_0_527[15:8]    = Image[626];
    assign  image_0_527[7:0]     = Image[627];

    assign  image_0_528[71:64]   = Image[562];
    assign  image_0_528[63:56]   = Image[563];
    assign  image_0_528[55:48]   = Image[564];
    assign  image_0_528[47:40]   = Image[594];
    assign  image_0_528[39:32]   = Image[595];
    assign  image_0_528[31:24]   = Image[596];
    assign  image_0_528[23:16]   = Image[626];
    assign  image_0_528[15:8]    = Image[627];
    assign  image_0_528[7:0]     = Image[628];

    assign  image_0_529[71:64]   = Image[563];
    assign  image_0_529[63:56]   = Image[564];
    assign  image_0_529[55:48]   = Image[565];
    assign  image_0_529[47:40]   = Image[595];
    assign  image_0_529[39:32]   = Image[596];
    assign  image_0_529[31:24]   = Image[597];
    assign  image_0_529[23:16]   = Image[627];
    assign  image_0_529[15:8]    = Image[628];
    assign  image_0_529[7:0]     = Image[629];

    assign  image_0_530[71:64]   = Image[564];
    assign  image_0_530[63:56]   = Image[565];
    assign  image_0_530[55:48]   = Image[566];
    assign  image_0_530[47:40]   = Image[596];
    assign  image_0_530[39:32]   = Image[597];
    assign  image_0_530[31:24]   = Image[598];
    assign  image_0_530[23:16]   = Image[628];
    assign  image_0_530[15:8]    = Image[629];
    assign  image_0_530[7:0]     = Image[630];

    assign  image_0_531[71:64]   = Image[565];
    assign  image_0_531[63:56]   = Image[566];
    assign  image_0_531[55:48]   = Image[567];
    assign  image_0_531[47:40]   = Image[597];
    assign  image_0_531[39:32]   = Image[598];
    assign  image_0_531[31:24]   = Image[599];
    assign  image_0_531[23:16]   = Image[629];
    assign  image_0_531[15:8]    = Image[630];
    assign  image_0_531[7:0]     = Image[631];

    assign  image_0_532[71:64]   = Image[566];
    assign  image_0_532[63:56]   = Image[567];
    assign  image_0_532[55:48]   = Image[568];
    assign  image_0_532[47:40]   = Image[598];
    assign  image_0_532[39:32]   = Image[599];
    assign  image_0_532[31:24]   = Image[600];
    assign  image_0_532[23:16]   = Image[630];
    assign  image_0_532[15:8]    = Image[631];
    assign  image_0_532[7:0]     = Image[632];

    assign  image_0_533[71:64]   = Image[567];
    assign  image_0_533[63:56]   = Image[568];
    assign  image_0_533[55:48]   = Image[569];
    assign  image_0_533[47:40]   = Image[599];
    assign  image_0_533[39:32]   = Image[600];
    assign  image_0_533[31:24]   = Image[601];
    assign  image_0_533[23:16]   = Image[631];
    assign  image_0_533[15:8]    = Image[632];
    assign  image_0_533[7:0]     = Image[633];

    assign  image_0_534[71:64]   = Image[568];
    assign  image_0_534[63:56]   = Image[569];
    assign  image_0_534[55:48]   = Image[570];
    assign  image_0_534[47:40]   = Image[600];
    assign  image_0_534[39:32]   = Image[601];
    assign  image_0_534[31:24]   = Image[602];
    assign  image_0_534[23:16]   = Image[632];
    assign  image_0_534[15:8]    = Image[633];
    assign  image_0_534[7:0]     = Image[634];

    assign  image_0_535[71:64]   = Image[569];
    assign  image_0_535[63:56]   = Image[570];
    assign  image_0_535[55:48]   = Image[571];
    assign  image_0_535[47:40]   = Image[601];
    assign  image_0_535[39:32]   = Image[602];
    assign  image_0_535[31:24]   = Image[603];
    assign  image_0_535[23:16]   = Image[633];
    assign  image_0_535[15:8]    = Image[634];
    assign  image_0_535[7:0]     = Image[635];

    assign  image_0_536[71:64]   = Image[570];
    assign  image_0_536[63:56]   = Image[571];
    assign  image_0_536[55:48]   = Image[572];
    assign  image_0_536[47:40]   = Image[602];
    assign  image_0_536[39:32]   = Image[603];
    assign  image_0_536[31:24]   = Image[604];
    assign  image_0_536[23:16]   = Image[634];
    assign  image_0_536[15:8]    = Image[635];
    assign  image_0_536[7:0]     = Image[636];

    assign  image_0_537[71:64]   = Image[571];
    assign  image_0_537[63:56]   = Image[572];
    assign  image_0_537[55:48]   = Image[573];
    assign  image_0_537[47:40]   = Image[603];
    assign  image_0_537[39:32]   = Image[604];
    assign  image_0_537[31:24]   = Image[605];
    assign  image_0_537[23:16]   = Image[635];
    assign  image_0_537[15:8]    = Image[636];
    assign  image_0_537[7:0]     = Image[637];

    assign  image_0_538[71:64]   = Image[572];
    assign  image_0_538[63:56]   = Image[573];
    assign  image_0_538[55:48]   = Image[574];
    assign  image_0_538[47:40]   = Image[604];
    assign  image_0_538[39:32]   = Image[605];
    assign  image_0_538[31:24]   = Image[606];
    assign  image_0_538[23:16]   = Image[636];
    assign  image_0_538[15:8]    = Image[637];
    assign  image_0_538[7:0]     = Image[638];

    assign  image_0_539[71:64]   = Image[573];
    assign  image_0_539[63:56]   = Image[574];
    assign  image_0_539[55:48]   = Image[575];
    assign  image_0_539[47:40]   = Image[605];
    assign  image_0_539[39:32]   = Image[606];
    assign  image_0_539[31:24]   = Image[607];
    assign  image_0_539[23:16]   = Image[637];
    assign  image_0_539[15:8]    = Image[638];
    assign  image_0_539[7:0]     = Image[639];

    assign  image_0_540[71:64]   = Image[576];
    assign  image_0_540[63:56]   = Image[577];
    assign  image_0_540[55:48]   = Image[578];
    assign  image_0_540[47:40]   = Image[608];
    assign  image_0_540[39:32]   = Image[609];
    assign  image_0_540[31:24]   = Image[610];
    assign  image_0_540[23:16]   = Image[640];
    assign  image_0_540[15:8]    = Image[641];
    assign  image_0_540[7:0]     = Image[642];

    assign  image_0_541[71:64]   = Image[577];
    assign  image_0_541[63:56]   = Image[578];
    assign  image_0_541[55:48]   = Image[579];
    assign  image_0_541[47:40]   = Image[609];
    assign  image_0_541[39:32]   = Image[610];
    assign  image_0_541[31:24]   = Image[611];
    assign  image_0_541[23:16]   = Image[641];
    assign  image_0_541[15:8]    = Image[642];
    assign  image_0_541[7:0]     = Image[643];

    assign  image_0_542[71:64]   = Image[578];
    assign  image_0_542[63:56]   = Image[579];
    assign  image_0_542[55:48]   = Image[580];
    assign  image_0_542[47:40]   = Image[610];
    assign  image_0_542[39:32]   = Image[611];
    assign  image_0_542[31:24]   = Image[612];
    assign  image_0_542[23:16]   = Image[642];
    assign  image_0_542[15:8]    = Image[643];
    assign  image_0_542[7:0]     = Image[644];

    assign  image_0_543[71:64]   = Image[579];
    assign  image_0_543[63:56]   = Image[580];
    assign  image_0_543[55:48]   = Image[581];
    assign  image_0_543[47:40]   = Image[611];
    assign  image_0_543[39:32]   = Image[612];
    assign  image_0_543[31:24]   = Image[613];
    assign  image_0_543[23:16]   = Image[643];
    assign  image_0_543[15:8]    = Image[644];
    assign  image_0_543[7:0]     = Image[645];

    assign  image_0_544[71:64]   = Image[580];
    assign  image_0_544[63:56]   = Image[581];
    assign  image_0_544[55:48]   = Image[582];
    assign  image_0_544[47:40]   = Image[612];
    assign  image_0_544[39:32]   = Image[613];
    assign  image_0_544[31:24]   = Image[614];
    assign  image_0_544[23:16]   = Image[644];
    assign  image_0_544[15:8]    = Image[645];
    assign  image_0_544[7:0]     = Image[646];

    assign  image_0_545[71:64]   = Image[581];
    assign  image_0_545[63:56]   = Image[582];
    assign  image_0_545[55:48]   = Image[583];
    assign  image_0_545[47:40]   = Image[613];
    assign  image_0_545[39:32]   = Image[614];
    assign  image_0_545[31:24]   = Image[615];
    assign  image_0_545[23:16]   = Image[645];
    assign  image_0_545[15:8]    = Image[646];
    assign  image_0_545[7:0]     = Image[647];

    assign  image_0_546[71:64]   = Image[582];
    assign  image_0_546[63:56]   = Image[583];
    assign  image_0_546[55:48]   = Image[584];
    assign  image_0_546[47:40]   = Image[614];
    assign  image_0_546[39:32]   = Image[615];
    assign  image_0_546[31:24]   = Image[616];
    assign  image_0_546[23:16]   = Image[646];
    assign  image_0_546[15:8]    = Image[647];
    assign  image_0_546[7:0]     = Image[648];

    assign  image_0_547[71:64]   = Image[583];
    assign  image_0_547[63:56]   = Image[584];
    assign  image_0_547[55:48]   = Image[585];
    assign  image_0_547[47:40]   = Image[615];
    assign  image_0_547[39:32]   = Image[616];
    assign  image_0_547[31:24]   = Image[617];
    assign  image_0_547[23:16]   = Image[647];
    assign  image_0_547[15:8]    = Image[648];
    assign  image_0_547[7:0]     = Image[649];

    assign  image_0_548[71:64]   = Image[584];
    assign  image_0_548[63:56]   = Image[585];
    assign  image_0_548[55:48]   = Image[586];
    assign  image_0_548[47:40]   = Image[616];
    assign  image_0_548[39:32]   = Image[617];
    assign  image_0_548[31:24]   = Image[618];
    assign  image_0_548[23:16]   = Image[648];
    assign  image_0_548[15:8]    = Image[649];
    assign  image_0_548[7:0]     = Image[650];

    assign  image_0_549[71:64]   = Image[585];
    assign  image_0_549[63:56]   = Image[586];
    assign  image_0_549[55:48]   = Image[587];
    assign  image_0_549[47:40]   = Image[617];
    assign  image_0_549[39:32]   = Image[618];
    assign  image_0_549[31:24]   = Image[619];
    assign  image_0_549[23:16]   = Image[649];
    assign  image_0_549[15:8]    = Image[650];
    assign  image_0_549[7:0]     = Image[651];

    assign  image_0_550[71:64]   = Image[586];
    assign  image_0_550[63:56]   = Image[587];
    assign  image_0_550[55:48]   = Image[588];
    assign  image_0_550[47:40]   = Image[618];
    assign  image_0_550[39:32]   = Image[619];
    assign  image_0_550[31:24]   = Image[620];
    assign  image_0_550[23:16]   = Image[650];
    assign  image_0_550[15:8]    = Image[651];
    assign  image_0_550[7:0]     = Image[652];

    assign  image_0_551[71:64]   = Image[587];
    assign  image_0_551[63:56]   = Image[588];
    assign  image_0_551[55:48]   = Image[589];
    assign  image_0_551[47:40]   = Image[619];
    assign  image_0_551[39:32]   = Image[620];
    assign  image_0_551[31:24]   = Image[621];
    assign  image_0_551[23:16]   = Image[651];
    assign  image_0_551[15:8]    = Image[652];
    assign  image_0_551[7:0]     = Image[653];

    assign  image_0_552[71:64]   = Image[588];
    assign  image_0_552[63:56]   = Image[589];
    assign  image_0_552[55:48]   = Image[590];
    assign  image_0_552[47:40]   = Image[620];
    assign  image_0_552[39:32]   = Image[621];
    assign  image_0_552[31:24]   = Image[622];
    assign  image_0_552[23:16]   = Image[652];
    assign  image_0_552[15:8]    = Image[653];
    assign  image_0_552[7:0]     = Image[654];

    assign  image_0_553[71:64]   = Image[589];
    assign  image_0_553[63:56]   = Image[590];
    assign  image_0_553[55:48]   = Image[591];
    assign  image_0_553[47:40]   = Image[621];
    assign  image_0_553[39:32]   = Image[622];
    assign  image_0_553[31:24]   = Image[623];
    assign  image_0_553[23:16]   = Image[653];
    assign  image_0_553[15:8]    = Image[654];
    assign  image_0_553[7:0]     = Image[655];

    assign  image_0_554[71:64]   = Image[590];
    assign  image_0_554[63:56]   = Image[591];
    assign  image_0_554[55:48]   = Image[592];
    assign  image_0_554[47:40]   = Image[622];
    assign  image_0_554[39:32]   = Image[623];
    assign  image_0_554[31:24]   = Image[624];
    assign  image_0_554[23:16]   = Image[654];
    assign  image_0_554[15:8]    = Image[655];
    assign  image_0_554[7:0]     = Image[656];

    assign  image_0_555[71:64]   = Image[591];
    assign  image_0_555[63:56]   = Image[592];
    assign  image_0_555[55:48]   = Image[593];
    assign  image_0_555[47:40]   = Image[623];
    assign  image_0_555[39:32]   = Image[624];
    assign  image_0_555[31:24]   = Image[625];
    assign  image_0_555[23:16]   = Image[655];
    assign  image_0_555[15:8]    = Image[656];
    assign  image_0_555[7:0]     = Image[657];

    assign  image_0_556[71:64]   = Image[592];
    assign  image_0_556[63:56]   = Image[593];
    assign  image_0_556[55:48]   = Image[594];
    assign  image_0_556[47:40]   = Image[624];
    assign  image_0_556[39:32]   = Image[625];
    assign  image_0_556[31:24]   = Image[626];
    assign  image_0_556[23:16]   = Image[656];
    assign  image_0_556[15:8]    = Image[657];
    assign  image_0_556[7:0]     = Image[658];

    assign  image_0_557[71:64]   = Image[593];
    assign  image_0_557[63:56]   = Image[594];
    assign  image_0_557[55:48]   = Image[595];
    assign  image_0_557[47:40]   = Image[625];
    assign  image_0_557[39:32]   = Image[626];
    assign  image_0_557[31:24]   = Image[627];
    assign  image_0_557[23:16]   = Image[657];
    assign  image_0_557[15:8]    = Image[658];
    assign  image_0_557[7:0]     = Image[659];

    assign  image_0_558[71:64]   = Image[594];
    assign  image_0_558[63:56]   = Image[595];
    assign  image_0_558[55:48]   = Image[596];
    assign  image_0_558[47:40]   = Image[626];
    assign  image_0_558[39:32]   = Image[627];
    assign  image_0_558[31:24]   = Image[628];
    assign  image_0_558[23:16]   = Image[658];
    assign  image_0_558[15:8]    = Image[659];
    assign  image_0_558[7:0]     = Image[660];

    assign  image_0_559[71:64]   = Image[595];
    assign  image_0_559[63:56]   = Image[596];
    assign  image_0_559[55:48]   = Image[597];
    assign  image_0_559[47:40]   = Image[627];
    assign  image_0_559[39:32]   = Image[628];
    assign  image_0_559[31:24]   = Image[629];
    assign  image_0_559[23:16]   = Image[659];
    assign  image_0_559[15:8]    = Image[660];
    assign  image_0_559[7:0]     = Image[661];

    assign  image_0_560[71:64]   = Image[596];
    assign  image_0_560[63:56]   = Image[597];
    assign  image_0_560[55:48]   = Image[598];
    assign  image_0_560[47:40]   = Image[628];
    assign  image_0_560[39:32]   = Image[629];
    assign  image_0_560[31:24]   = Image[630];
    assign  image_0_560[23:16]   = Image[660];
    assign  image_0_560[15:8]    = Image[661];
    assign  image_0_560[7:0]     = Image[662];

    assign  image_0_561[71:64]   = Image[597];
    assign  image_0_561[63:56]   = Image[598];
    assign  image_0_561[55:48]   = Image[599];
    assign  image_0_561[47:40]   = Image[629];
    assign  image_0_561[39:32]   = Image[630];
    assign  image_0_561[31:24]   = Image[631];
    assign  image_0_561[23:16]   = Image[661];
    assign  image_0_561[15:8]    = Image[662];
    assign  image_0_561[7:0]     = Image[663];

    assign  image_0_562[71:64]   = Image[598];
    assign  image_0_562[63:56]   = Image[599];
    assign  image_0_562[55:48]   = Image[600];
    assign  image_0_562[47:40]   = Image[630];
    assign  image_0_562[39:32]   = Image[631];
    assign  image_0_562[31:24]   = Image[632];
    assign  image_0_562[23:16]   = Image[662];
    assign  image_0_562[15:8]    = Image[663];
    assign  image_0_562[7:0]     = Image[664];

    assign  image_0_563[71:64]   = Image[599];
    assign  image_0_563[63:56]   = Image[600];
    assign  image_0_563[55:48]   = Image[601];
    assign  image_0_563[47:40]   = Image[631];
    assign  image_0_563[39:32]   = Image[632];
    assign  image_0_563[31:24]   = Image[633];
    assign  image_0_563[23:16]   = Image[663];
    assign  image_0_563[15:8]    = Image[664];
    assign  image_0_563[7:0]     = Image[665];

    assign  image_0_564[71:64]   = Image[600];
    assign  image_0_564[63:56]   = Image[601];
    assign  image_0_564[55:48]   = Image[602];
    assign  image_0_564[47:40]   = Image[632];
    assign  image_0_564[39:32]   = Image[633];
    assign  image_0_564[31:24]   = Image[634];
    assign  image_0_564[23:16]   = Image[664];
    assign  image_0_564[15:8]    = Image[665];
    assign  image_0_564[7:0]     = Image[666];

    assign  image_0_565[71:64]   = Image[601];
    assign  image_0_565[63:56]   = Image[602];
    assign  image_0_565[55:48]   = Image[603];
    assign  image_0_565[47:40]   = Image[633];
    assign  image_0_565[39:32]   = Image[634];
    assign  image_0_565[31:24]   = Image[635];
    assign  image_0_565[23:16]   = Image[665];
    assign  image_0_565[15:8]    = Image[666];
    assign  image_0_565[7:0]     = Image[667];

    assign  image_0_566[71:64]   = Image[602];
    assign  image_0_566[63:56]   = Image[603];
    assign  image_0_566[55:48]   = Image[604];
    assign  image_0_566[47:40]   = Image[634];
    assign  image_0_566[39:32]   = Image[635];
    assign  image_0_566[31:24]   = Image[636];
    assign  image_0_566[23:16]   = Image[666];
    assign  image_0_566[15:8]    = Image[667];
    assign  image_0_566[7:0]     = Image[668];

    assign  image_0_567[71:64]   = Image[603];
    assign  image_0_567[63:56]   = Image[604];
    assign  image_0_567[55:48]   = Image[605];
    assign  image_0_567[47:40]   = Image[635];
    assign  image_0_567[39:32]   = Image[636];
    assign  image_0_567[31:24]   = Image[637];
    assign  image_0_567[23:16]   = Image[667];
    assign  image_0_567[15:8]    = Image[668];
    assign  image_0_567[7:0]     = Image[669];

    assign  image_0_568[71:64]   = Image[604];
    assign  image_0_568[63:56]   = Image[605];
    assign  image_0_568[55:48]   = Image[606];
    assign  image_0_568[47:40]   = Image[636];
    assign  image_0_568[39:32]   = Image[637];
    assign  image_0_568[31:24]   = Image[638];
    assign  image_0_568[23:16]   = Image[668];
    assign  image_0_568[15:8]    = Image[669];
    assign  image_0_568[7:0]     = Image[670];

    assign  image_0_569[71:64]   = Image[605];
    assign  image_0_569[63:56]   = Image[606];
    assign  image_0_569[55:48]   = Image[607];
    assign  image_0_569[47:40]   = Image[637];
    assign  image_0_569[39:32]   = Image[638];
    assign  image_0_569[31:24]   = Image[639];
    assign  image_0_569[23:16]   = Image[669];
    assign  image_0_569[15:8]    = Image[670];
    assign  image_0_569[7:0]     = Image[671];

    assign  image_0_570[71:64]   = Image[608];
    assign  image_0_570[63:56]   = Image[609];
    assign  image_0_570[55:48]   = Image[610];
    assign  image_0_570[47:40]   = Image[640];
    assign  image_0_570[39:32]   = Image[641];
    assign  image_0_570[31:24]   = Image[642];
    assign  image_0_570[23:16]   = Image[672];
    assign  image_0_570[15:8]    = Image[673];
    assign  image_0_570[7:0]     = Image[674];

    assign  image_0_571[71:64]   = Image[609];
    assign  image_0_571[63:56]   = Image[610];
    assign  image_0_571[55:48]   = Image[611];
    assign  image_0_571[47:40]   = Image[641];
    assign  image_0_571[39:32]   = Image[642];
    assign  image_0_571[31:24]   = Image[643];
    assign  image_0_571[23:16]   = Image[673];
    assign  image_0_571[15:8]    = Image[674];
    assign  image_0_571[7:0]     = Image[675];

    assign  image_0_572[71:64]   = Image[610];
    assign  image_0_572[63:56]   = Image[611];
    assign  image_0_572[55:48]   = Image[612];
    assign  image_0_572[47:40]   = Image[642];
    assign  image_0_572[39:32]   = Image[643];
    assign  image_0_572[31:24]   = Image[644];
    assign  image_0_572[23:16]   = Image[674];
    assign  image_0_572[15:8]    = Image[675];
    assign  image_0_572[7:0]     = Image[676];

    assign  image_0_573[71:64]   = Image[611];
    assign  image_0_573[63:56]   = Image[612];
    assign  image_0_573[55:48]   = Image[613];
    assign  image_0_573[47:40]   = Image[643];
    assign  image_0_573[39:32]   = Image[644];
    assign  image_0_573[31:24]   = Image[645];
    assign  image_0_573[23:16]   = Image[675];
    assign  image_0_573[15:8]    = Image[676];
    assign  image_0_573[7:0]     = Image[677];

    assign  image_0_574[71:64]   = Image[612];
    assign  image_0_574[63:56]   = Image[613];
    assign  image_0_574[55:48]   = Image[614];
    assign  image_0_574[47:40]   = Image[644];
    assign  image_0_574[39:32]   = Image[645];
    assign  image_0_574[31:24]   = Image[646];
    assign  image_0_574[23:16]   = Image[676];
    assign  image_0_574[15:8]    = Image[677];
    assign  image_0_574[7:0]     = Image[678];

    assign  image_0_575[71:64]   = Image[613];
    assign  image_0_575[63:56]   = Image[614];
    assign  image_0_575[55:48]   = Image[615];
    assign  image_0_575[47:40]   = Image[645];
    assign  image_0_575[39:32]   = Image[646];
    assign  image_0_575[31:24]   = Image[647];
    assign  image_0_575[23:16]   = Image[677];
    assign  image_0_575[15:8]    = Image[678];
    assign  image_0_575[7:0]     = Image[679];

    assign  image_0_576[71:64]   = Image[614];
    assign  image_0_576[63:56]   = Image[615];
    assign  image_0_576[55:48]   = Image[616];
    assign  image_0_576[47:40]   = Image[646];
    assign  image_0_576[39:32]   = Image[647];
    assign  image_0_576[31:24]   = Image[648];
    assign  image_0_576[23:16]   = Image[678];
    assign  image_0_576[15:8]    = Image[679];
    assign  image_0_576[7:0]     = Image[680];

    assign  image_0_577[71:64]   = Image[615];
    assign  image_0_577[63:56]   = Image[616];
    assign  image_0_577[55:48]   = Image[617];
    assign  image_0_577[47:40]   = Image[647];
    assign  image_0_577[39:32]   = Image[648];
    assign  image_0_577[31:24]   = Image[649];
    assign  image_0_577[23:16]   = Image[679];
    assign  image_0_577[15:8]    = Image[680];
    assign  image_0_577[7:0]     = Image[681];

    assign  image_0_578[71:64]   = Image[616];
    assign  image_0_578[63:56]   = Image[617];
    assign  image_0_578[55:48]   = Image[618];
    assign  image_0_578[47:40]   = Image[648];
    assign  image_0_578[39:32]   = Image[649];
    assign  image_0_578[31:24]   = Image[650];
    assign  image_0_578[23:16]   = Image[680];
    assign  image_0_578[15:8]    = Image[681];
    assign  image_0_578[7:0]     = Image[682];

    assign  image_0_579[71:64]   = Image[617];
    assign  image_0_579[63:56]   = Image[618];
    assign  image_0_579[55:48]   = Image[619];
    assign  image_0_579[47:40]   = Image[649];
    assign  image_0_579[39:32]   = Image[650];
    assign  image_0_579[31:24]   = Image[651];
    assign  image_0_579[23:16]   = Image[681];
    assign  image_0_579[15:8]    = Image[682];
    assign  image_0_579[7:0]     = Image[683];

    assign  image_0_580[71:64]   = Image[618];
    assign  image_0_580[63:56]   = Image[619];
    assign  image_0_580[55:48]   = Image[620];
    assign  image_0_580[47:40]   = Image[650];
    assign  image_0_580[39:32]   = Image[651];
    assign  image_0_580[31:24]   = Image[652];
    assign  image_0_580[23:16]   = Image[682];
    assign  image_0_580[15:8]    = Image[683];
    assign  image_0_580[7:0]     = Image[684];

    assign  image_0_581[71:64]   = Image[619];
    assign  image_0_581[63:56]   = Image[620];
    assign  image_0_581[55:48]   = Image[621];
    assign  image_0_581[47:40]   = Image[651];
    assign  image_0_581[39:32]   = Image[652];
    assign  image_0_581[31:24]   = Image[653];
    assign  image_0_581[23:16]   = Image[683];
    assign  image_0_581[15:8]    = Image[684];
    assign  image_0_581[7:0]     = Image[685];

    assign  image_0_582[71:64]   = Image[620];
    assign  image_0_582[63:56]   = Image[621];
    assign  image_0_582[55:48]   = Image[622];
    assign  image_0_582[47:40]   = Image[652];
    assign  image_0_582[39:32]   = Image[653];
    assign  image_0_582[31:24]   = Image[654];
    assign  image_0_582[23:16]   = Image[684];
    assign  image_0_582[15:8]    = Image[685];
    assign  image_0_582[7:0]     = Image[686];

    assign  image_0_583[71:64]   = Image[621];
    assign  image_0_583[63:56]   = Image[622];
    assign  image_0_583[55:48]   = Image[623];
    assign  image_0_583[47:40]   = Image[653];
    assign  image_0_583[39:32]   = Image[654];
    assign  image_0_583[31:24]   = Image[655];
    assign  image_0_583[23:16]   = Image[685];
    assign  image_0_583[15:8]    = Image[686];
    assign  image_0_583[7:0]     = Image[687];

    assign  image_0_584[71:64]   = Image[622];
    assign  image_0_584[63:56]   = Image[623];
    assign  image_0_584[55:48]   = Image[624];
    assign  image_0_584[47:40]   = Image[654];
    assign  image_0_584[39:32]   = Image[655];
    assign  image_0_584[31:24]   = Image[656];
    assign  image_0_584[23:16]   = Image[686];
    assign  image_0_584[15:8]    = Image[687];
    assign  image_0_584[7:0]     = Image[688];

    assign  image_0_585[71:64]   = Image[623];
    assign  image_0_585[63:56]   = Image[624];
    assign  image_0_585[55:48]   = Image[625];
    assign  image_0_585[47:40]   = Image[655];
    assign  image_0_585[39:32]   = Image[656];
    assign  image_0_585[31:24]   = Image[657];
    assign  image_0_585[23:16]   = Image[687];
    assign  image_0_585[15:8]    = Image[688];
    assign  image_0_585[7:0]     = Image[689];

    assign  image_0_586[71:64]   = Image[624];
    assign  image_0_586[63:56]   = Image[625];
    assign  image_0_586[55:48]   = Image[626];
    assign  image_0_586[47:40]   = Image[656];
    assign  image_0_586[39:32]   = Image[657];
    assign  image_0_586[31:24]   = Image[658];
    assign  image_0_586[23:16]   = Image[688];
    assign  image_0_586[15:8]    = Image[689];
    assign  image_0_586[7:0]     = Image[690];

    assign  image_0_587[71:64]   = Image[625];
    assign  image_0_587[63:56]   = Image[626];
    assign  image_0_587[55:48]   = Image[627];
    assign  image_0_587[47:40]   = Image[657];
    assign  image_0_587[39:32]   = Image[658];
    assign  image_0_587[31:24]   = Image[659];
    assign  image_0_587[23:16]   = Image[689];
    assign  image_0_587[15:8]    = Image[690];
    assign  image_0_587[7:0]     = Image[691];

    assign  image_0_588[71:64]   = Image[626];
    assign  image_0_588[63:56]   = Image[627];
    assign  image_0_588[55:48]   = Image[628];
    assign  image_0_588[47:40]   = Image[658];
    assign  image_0_588[39:32]   = Image[659];
    assign  image_0_588[31:24]   = Image[660];
    assign  image_0_588[23:16]   = Image[690];
    assign  image_0_588[15:8]    = Image[691];
    assign  image_0_588[7:0]     = Image[692];

    assign  image_0_589[71:64]   = Image[627];
    assign  image_0_589[63:56]   = Image[628];
    assign  image_0_589[55:48]   = Image[629];
    assign  image_0_589[47:40]   = Image[659];
    assign  image_0_589[39:32]   = Image[660];
    assign  image_0_589[31:24]   = Image[661];
    assign  image_0_589[23:16]   = Image[691];
    assign  image_0_589[15:8]    = Image[692];
    assign  image_0_589[7:0]     = Image[693];

    assign  image_0_590[71:64]   = Image[628];
    assign  image_0_590[63:56]   = Image[629];
    assign  image_0_590[55:48]   = Image[630];
    assign  image_0_590[47:40]   = Image[660];
    assign  image_0_590[39:32]   = Image[661];
    assign  image_0_590[31:24]   = Image[662];
    assign  image_0_590[23:16]   = Image[692];
    assign  image_0_590[15:8]    = Image[693];
    assign  image_0_590[7:0]     = Image[694];

    assign  image_0_591[71:64]   = Image[629];
    assign  image_0_591[63:56]   = Image[630];
    assign  image_0_591[55:48]   = Image[631];
    assign  image_0_591[47:40]   = Image[661];
    assign  image_0_591[39:32]   = Image[662];
    assign  image_0_591[31:24]   = Image[663];
    assign  image_0_591[23:16]   = Image[693];
    assign  image_0_591[15:8]    = Image[694];
    assign  image_0_591[7:0]     = Image[695];

    assign  image_0_592[71:64]   = Image[630];
    assign  image_0_592[63:56]   = Image[631];
    assign  image_0_592[55:48]   = Image[632];
    assign  image_0_592[47:40]   = Image[662];
    assign  image_0_592[39:32]   = Image[663];
    assign  image_0_592[31:24]   = Image[664];
    assign  image_0_592[23:16]   = Image[694];
    assign  image_0_592[15:8]    = Image[695];
    assign  image_0_592[7:0]     = Image[696];

    assign  image_0_593[71:64]   = Image[631];
    assign  image_0_593[63:56]   = Image[632];
    assign  image_0_593[55:48]   = Image[633];
    assign  image_0_593[47:40]   = Image[663];
    assign  image_0_593[39:32]   = Image[664];
    assign  image_0_593[31:24]   = Image[665];
    assign  image_0_593[23:16]   = Image[695];
    assign  image_0_593[15:8]    = Image[696];
    assign  image_0_593[7:0]     = Image[697];

    assign  image_0_594[71:64]   = Image[632];
    assign  image_0_594[63:56]   = Image[633];
    assign  image_0_594[55:48]   = Image[634];
    assign  image_0_594[47:40]   = Image[664];
    assign  image_0_594[39:32]   = Image[665];
    assign  image_0_594[31:24]   = Image[666];
    assign  image_0_594[23:16]   = Image[696];
    assign  image_0_594[15:8]    = Image[697];
    assign  image_0_594[7:0]     = Image[698];

    assign  image_0_595[71:64]   = Image[633];
    assign  image_0_595[63:56]   = Image[634];
    assign  image_0_595[55:48]   = Image[635];
    assign  image_0_595[47:40]   = Image[665];
    assign  image_0_595[39:32]   = Image[666];
    assign  image_0_595[31:24]   = Image[667];
    assign  image_0_595[23:16]   = Image[697];
    assign  image_0_595[15:8]    = Image[698];
    assign  image_0_595[7:0]     = Image[699];

    assign  image_0_596[71:64]   = Image[634];
    assign  image_0_596[63:56]   = Image[635];
    assign  image_0_596[55:48]   = Image[636];
    assign  image_0_596[47:40]   = Image[666];
    assign  image_0_596[39:32]   = Image[667];
    assign  image_0_596[31:24]   = Image[668];
    assign  image_0_596[23:16]   = Image[698];
    assign  image_0_596[15:8]    = Image[699];
    assign  image_0_596[7:0]     = Image[700];

    assign  image_0_597[71:64]   = Image[635];
    assign  image_0_597[63:56]   = Image[636];
    assign  image_0_597[55:48]   = Image[637];
    assign  image_0_597[47:40]   = Image[667];
    assign  image_0_597[39:32]   = Image[668];
    assign  image_0_597[31:24]   = Image[669];
    assign  image_0_597[23:16]   = Image[699];
    assign  image_0_597[15:8]    = Image[700];
    assign  image_0_597[7:0]     = Image[701];

    assign  image_0_598[71:64]   = Image[636];
    assign  image_0_598[63:56]   = Image[637];
    assign  image_0_598[55:48]   = Image[638];
    assign  image_0_598[47:40]   = Image[668];
    assign  image_0_598[39:32]   = Image[669];
    assign  image_0_598[31:24]   = Image[670];
    assign  image_0_598[23:16]   = Image[700];
    assign  image_0_598[15:8]    = Image[701];
    assign  image_0_598[7:0]     = Image[702];

    assign  image_0_599[71:64]   = Image[637];
    assign  image_0_599[63:56]   = Image[638];
    assign  image_0_599[55:48]   = Image[639];
    assign  image_0_599[47:40]   = Image[669];
    assign  image_0_599[39:32]   = Image[670];
    assign  image_0_599[31:24]   = Image[671];
    assign  image_0_599[23:16]   = Image[701];
    assign  image_0_599[15:8]    = Image[702];
    assign  image_0_599[7:0]     = Image[703];

    assign  image_0_600[71:64]   = Image[640];
    assign  image_0_600[63:56]   = Image[641];
    assign  image_0_600[55:48]   = Image[642];
    assign  image_0_600[47:40]   = Image[672];
    assign  image_0_600[39:32]   = Image[673];
    assign  image_0_600[31:24]   = Image[674];
    assign  image_0_600[23:16]   = Image[704];
    assign  image_0_600[15:8]    = Image[705];
    assign  image_0_600[7:0]     = Image[706];

    assign  image_0_601[71:64]   = Image[641];
    assign  image_0_601[63:56]   = Image[642];
    assign  image_0_601[55:48]   = Image[643];
    assign  image_0_601[47:40]   = Image[673];
    assign  image_0_601[39:32]   = Image[674];
    assign  image_0_601[31:24]   = Image[675];
    assign  image_0_601[23:16]   = Image[705];
    assign  image_0_601[15:8]    = Image[706];
    assign  image_0_601[7:0]     = Image[707];

    assign  image_0_602[71:64]   = Image[642];
    assign  image_0_602[63:56]   = Image[643];
    assign  image_0_602[55:48]   = Image[644];
    assign  image_0_602[47:40]   = Image[674];
    assign  image_0_602[39:32]   = Image[675];
    assign  image_0_602[31:24]   = Image[676];
    assign  image_0_602[23:16]   = Image[706];
    assign  image_0_602[15:8]    = Image[707];
    assign  image_0_602[7:0]     = Image[708];

    assign  image_0_603[71:64]   = Image[643];
    assign  image_0_603[63:56]   = Image[644];
    assign  image_0_603[55:48]   = Image[645];
    assign  image_0_603[47:40]   = Image[675];
    assign  image_0_603[39:32]   = Image[676];
    assign  image_0_603[31:24]   = Image[677];
    assign  image_0_603[23:16]   = Image[707];
    assign  image_0_603[15:8]    = Image[708];
    assign  image_0_603[7:0]     = Image[709];

    assign  image_0_604[71:64]   = Image[644];
    assign  image_0_604[63:56]   = Image[645];
    assign  image_0_604[55:48]   = Image[646];
    assign  image_0_604[47:40]   = Image[676];
    assign  image_0_604[39:32]   = Image[677];
    assign  image_0_604[31:24]   = Image[678];
    assign  image_0_604[23:16]   = Image[708];
    assign  image_0_604[15:8]    = Image[709];
    assign  image_0_604[7:0]     = Image[710];

    assign  image_0_605[71:64]   = Image[645];
    assign  image_0_605[63:56]   = Image[646];
    assign  image_0_605[55:48]   = Image[647];
    assign  image_0_605[47:40]   = Image[677];
    assign  image_0_605[39:32]   = Image[678];
    assign  image_0_605[31:24]   = Image[679];
    assign  image_0_605[23:16]   = Image[709];
    assign  image_0_605[15:8]    = Image[710];
    assign  image_0_605[7:0]     = Image[711];

    assign  image_0_606[71:64]   = Image[646];
    assign  image_0_606[63:56]   = Image[647];
    assign  image_0_606[55:48]   = Image[648];
    assign  image_0_606[47:40]   = Image[678];
    assign  image_0_606[39:32]   = Image[679];
    assign  image_0_606[31:24]   = Image[680];
    assign  image_0_606[23:16]   = Image[710];
    assign  image_0_606[15:8]    = Image[711];
    assign  image_0_606[7:0]     = Image[712];

    assign  image_0_607[71:64]   = Image[647];
    assign  image_0_607[63:56]   = Image[648];
    assign  image_0_607[55:48]   = Image[649];
    assign  image_0_607[47:40]   = Image[679];
    assign  image_0_607[39:32]   = Image[680];
    assign  image_0_607[31:24]   = Image[681];
    assign  image_0_607[23:16]   = Image[711];
    assign  image_0_607[15:8]    = Image[712];
    assign  image_0_607[7:0]     = Image[713];

    assign  image_0_608[71:64]   = Image[648];
    assign  image_0_608[63:56]   = Image[649];
    assign  image_0_608[55:48]   = Image[650];
    assign  image_0_608[47:40]   = Image[680];
    assign  image_0_608[39:32]   = Image[681];
    assign  image_0_608[31:24]   = Image[682];
    assign  image_0_608[23:16]   = Image[712];
    assign  image_0_608[15:8]    = Image[713];
    assign  image_0_608[7:0]     = Image[714];

    assign  image_0_609[71:64]   = Image[649];
    assign  image_0_609[63:56]   = Image[650];
    assign  image_0_609[55:48]   = Image[651];
    assign  image_0_609[47:40]   = Image[681];
    assign  image_0_609[39:32]   = Image[682];
    assign  image_0_609[31:24]   = Image[683];
    assign  image_0_609[23:16]   = Image[713];
    assign  image_0_609[15:8]    = Image[714];
    assign  image_0_609[7:0]     = Image[715];

    assign  image_0_610[71:64]   = Image[650];
    assign  image_0_610[63:56]   = Image[651];
    assign  image_0_610[55:48]   = Image[652];
    assign  image_0_610[47:40]   = Image[682];
    assign  image_0_610[39:32]   = Image[683];
    assign  image_0_610[31:24]   = Image[684];
    assign  image_0_610[23:16]   = Image[714];
    assign  image_0_610[15:8]    = Image[715];
    assign  image_0_610[7:0]     = Image[716];

    assign  image_0_611[71:64]   = Image[651];
    assign  image_0_611[63:56]   = Image[652];
    assign  image_0_611[55:48]   = Image[653];
    assign  image_0_611[47:40]   = Image[683];
    assign  image_0_611[39:32]   = Image[684];
    assign  image_0_611[31:24]   = Image[685];
    assign  image_0_611[23:16]   = Image[715];
    assign  image_0_611[15:8]    = Image[716];
    assign  image_0_611[7:0]     = Image[717];

    assign  image_0_612[71:64]   = Image[652];
    assign  image_0_612[63:56]   = Image[653];
    assign  image_0_612[55:48]   = Image[654];
    assign  image_0_612[47:40]   = Image[684];
    assign  image_0_612[39:32]   = Image[685];
    assign  image_0_612[31:24]   = Image[686];
    assign  image_0_612[23:16]   = Image[716];
    assign  image_0_612[15:8]    = Image[717];
    assign  image_0_612[7:0]     = Image[718];

    assign  image_0_613[71:64]   = Image[653];
    assign  image_0_613[63:56]   = Image[654];
    assign  image_0_613[55:48]   = Image[655];
    assign  image_0_613[47:40]   = Image[685];
    assign  image_0_613[39:32]   = Image[686];
    assign  image_0_613[31:24]   = Image[687];
    assign  image_0_613[23:16]   = Image[717];
    assign  image_0_613[15:8]    = Image[718];
    assign  image_0_613[7:0]     = Image[719];

    assign  image_0_614[71:64]   = Image[654];
    assign  image_0_614[63:56]   = Image[655];
    assign  image_0_614[55:48]   = Image[656];
    assign  image_0_614[47:40]   = Image[686];
    assign  image_0_614[39:32]   = Image[687];
    assign  image_0_614[31:24]   = Image[688];
    assign  image_0_614[23:16]   = Image[718];
    assign  image_0_614[15:8]    = Image[719];
    assign  image_0_614[7:0]     = Image[720];

    assign  image_0_615[71:64]   = Image[655];
    assign  image_0_615[63:56]   = Image[656];
    assign  image_0_615[55:48]   = Image[657];
    assign  image_0_615[47:40]   = Image[687];
    assign  image_0_615[39:32]   = Image[688];
    assign  image_0_615[31:24]   = Image[689];
    assign  image_0_615[23:16]   = Image[719];
    assign  image_0_615[15:8]    = Image[720];
    assign  image_0_615[7:0]     = Image[721];

    assign  image_0_616[71:64]   = Image[656];
    assign  image_0_616[63:56]   = Image[657];
    assign  image_0_616[55:48]   = Image[658];
    assign  image_0_616[47:40]   = Image[688];
    assign  image_0_616[39:32]   = Image[689];
    assign  image_0_616[31:24]   = Image[690];
    assign  image_0_616[23:16]   = Image[720];
    assign  image_0_616[15:8]    = Image[721];
    assign  image_0_616[7:0]     = Image[722];

    assign  image_0_617[71:64]   = Image[657];
    assign  image_0_617[63:56]   = Image[658];
    assign  image_0_617[55:48]   = Image[659];
    assign  image_0_617[47:40]   = Image[689];
    assign  image_0_617[39:32]   = Image[690];
    assign  image_0_617[31:24]   = Image[691];
    assign  image_0_617[23:16]   = Image[721];
    assign  image_0_617[15:8]    = Image[722];
    assign  image_0_617[7:0]     = Image[723];

    assign  image_0_618[71:64]   = Image[658];
    assign  image_0_618[63:56]   = Image[659];
    assign  image_0_618[55:48]   = Image[660];
    assign  image_0_618[47:40]   = Image[690];
    assign  image_0_618[39:32]   = Image[691];
    assign  image_0_618[31:24]   = Image[692];
    assign  image_0_618[23:16]   = Image[722];
    assign  image_0_618[15:8]    = Image[723];
    assign  image_0_618[7:0]     = Image[724];

    assign  image_0_619[71:64]   = Image[659];
    assign  image_0_619[63:56]   = Image[660];
    assign  image_0_619[55:48]   = Image[661];
    assign  image_0_619[47:40]   = Image[691];
    assign  image_0_619[39:32]   = Image[692];
    assign  image_0_619[31:24]   = Image[693];
    assign  image_0_619[23:16]   = Image[723];
    assign  image_0_619[15:8]    = Image[724];
    assign  image_0_619[7:0]     = Image[725];

    assign  image_0_620[71:64]   = Image[660];
    assign  image_0_620[63:56]   = Image[661];
    assign  image_0_620[55:48]   = Image[662];
    assign  image_0_620[47:40]   = Image[692];
    assign  image_0_620[39:32]   = Image[693];
    assign  image_0_620[31:24]   = Image[694];
    assign  image_0_620[23:16]   = Image[724];
    assign  image_0_620[15:8]    = Image[725];
    assign  image_0_620[7:0]     = Image[726];

    assign  image_0_621[71:64]   = Image[661];
    assign  image_0_621[63:56]   = Image[662];
    assign  image_0_621[55:48]   = Image[663];
    assign  image_0_621[47:40]   = Image[693];
    assign  image_0_621[39:32]   = Image[694];
    assign  image_0_621[31:24]   = Image[695];
    assign  image_0_621[23:16]   = Image[725];
    assign  image_0_621[15:8]    = Image[726];
    assign  image_0_621[7:0]     = Image[727];

    assign  image_0_622[71:64]   = Image[662];
    assign  image_0_622[63:56]   = Image[663];
    assign  image_0_622[55:48]   = Image[664];
    assign  image_0_622[47:40]   = Image[694];
    assign  image_0_622[39:32]   = Image[695];
    assign  image_0_622[31:24]   = Image[696];
    assign  image_0_622[23:16]   = Image[726];
    assign  image_0_622[15:8]    = Image[727];
    assign  image_0_622[7:0]     = Image[728];

    assign  image_0_623[71:64]   = Image[663];
    assign  image_0_623[63:56]   = Image[664];
    assign  image_0_623[55:48]   = Image[665];
    assign  image_0_623[47:40]   = Image[695];
    assign  image_0_623[39:32]   = Image[696];
    assign  image_0_623[31:24]   = Image[697];
    assign  image_0_623[23:16]   = Image[727];
    assign  image_0_623[15:8]    = Image[728];
    assign  image_0_623[7:0]     = Image[729];

    assign  image_0_624[71:64]   = Image[664];
    assign  image_0_624[63:56]   = Image[665];
    assign  image_0_624[55:48]   = Image[666];
    assign  image_0_624[47:40]   = Image[696];
    assign  image_0_624[39:32]   = Image[697];
    assign  image_0_624[31:24]   = Image[698];
    assign  image_0_624[23:16]   = Image[728];
    assign  image_0_624[15:8]    = Image[729];
    assign  image_0_624[7:0]     = Image[730];

    assign  image_0_625[71:64]   = Image[665];
    assign  image_0_625[63:56]   = Image[666];
    assign  image_0_625[55:48]   = Image[667];
    assign  image_0_625[47:40]   = Image[697];
    assign  image_0_625[39:32]   = Image[698];
    assign  image_0_625[31:24]   = Image[699];
    assign  image_0_625[23:16]   = Image[729];
    assign  image_0_625[15:8]    = Image[730];
    assign  image_0_625[7:0]     = Image[731];

    assign  image_0_626[71:64]   = Image[666];
    assign  image_0_626[63:56]   = Image[667];
    assign  image_0_626[55:48]   = Image[668];
    assign  image_0_626[47:40]   = Image[698];
    assign  image_0_626[39:32]   = Image[699];
    assign  image_0_626[31:24]   = Image[700];
    assign  image_0_626[23:16]   = Image[730];
    assign  image_0_626[15:8]    = Image[731];
    assign  image_0_626[7:0]     = Image[732];

    assign  image_0_627[71:64]   = Image[667];
    assign  image_0_627[63:56]   = Image[668];
    assign  image_0_627[55:48]   = Image[669];
    assign  image_0_627[47:40]   = Image[699];
    assign  image_0_627[39:32]   = Image[700];
    assign  image_0_627[31:24]   = Image[701];
    assign  image_0_627[23:16]   = Image[731];
    assign  image_0_627[15:8]    = Image[732];
    assign  image_0_627[7:0]     = Image[733];

    assign  image_0_628[71:64]   = Image[668];
    assign  image_0_628[63:56]   = Image[669];
    assign  image_0_628[55:48]   = Image[670];
    assign  image_0_628[47:40]   = Image[700];
    assign  image_0_628[39:32]   = Image[701];
    assign  image_0_628[31:24]   = Image[702];
    assign  image_0_628[23:16]   = Image[732];
    assign  image_0_628[15:8]    = Image[733];
    assign  image_0_628[7:0]     = Image[734];

    assign  image_0_629[71:64]   = Image[669];
    assign  image_0_629[63:56]   = Image[670];
    assign  image_0_629[55:48]   = Image[671];
    assign  image_0_629[47:40]   = Image[701];
    assign  image_0_629[39:32]   = Image[702];
    assign  image_0_629[31:24]   = Image[703];
    assign  image_0_629[23:16]   = Image[733];
    assign  image_0_629[15:8]    = Image[734];
    assign  image_0_629[7:0]     = Image[735];

    assign  image_0_630[71:64]   = Image[672];
    assign  image_0_630[63:56]   = Image[673];
    assign  image_0_630[55:48]   = Image[674];
    assign  image_0_630[47:40]   = Image[704];
    assign  image_0_630[39:32]   = Image[705];
    assign  image_0_630[31:24]   = Image[706];
    assign  image_0_630[23:16]   = Image[736];
    assign  image_0_630[15:8]    = Image[737];
    assign  image_0_630[7:0]     = Image[738];

    assign  image_0_631[71:64]   = Image[673];
    assign  image_0_631[63:56]   = Image[674];
    assign  image_0_631[55:48]   = Image[675];
    assign  image_0_631[47:40]   = Image[705];
    assign  image_0_631[39:32]   = Image[706];
    assign  image_0_631[31:24]   = Image[707];
    assign  image_0_631[23:16]   = Image[737];
    assign  image_0_631[15:8]    = Image[738];
    assign  image_0_631[7:0]     = Image[739];

    assign  image_0_632[71:64]   = Image[674];
    assign  image_0_632[63:56]   = Image[675];
    assign  image_0_632[55:48]   = Image[676];
    assign  image_0_632[47:40]   = Image[706];
    assign  image_0_632[39:32]   = Image[707];
    assign  image_0_632[31:24]   = Image[708];
    assign  image_0_632[23:16]   = Image[738];
    assign  image_0_632[15:8]    = Image[739];
    assign  image_0_632[7:0]     = Image[740];

    assign  image_0_633[71:64]   = Image[675];
    assign  image_0_633[63:56]   = Image[676];
    assign  image_0_633[55:48]   = Image[677];
    assign  image_0_633[47:40]   = Image[707];
    assign  image_0_633[39:32]   = Image[708];
    assign  image_0_633[31:24]   = Image[709];
    assign  image_0_633[23:16]   = Image[739];
    assign  image_0_633[15:8]    = Image[740];
    assign  image_0_633[7:0]     = Image[741];

    assign  image_0_634[71:64]   = Image[676];
    assign  image_0_634[63:56]   = Image[677];
    assign  image_0_634[55:48]   = Image[678];
    assign  image_0_634[47:40]   = Image[708];
    assign  image_0_634[39:32]   = Image[709];
    assign  image_0_634[31:24]   = Image[710];
    assign  image_0_634[23:16]   = Image[740];
    assign  image_0_634[15:8]    = Image[741];
    assign  image_0_634[7:0]     = Image[742];

    assign  image_0_635[71:64]   = Image[677];
    assign  image_0_635[63:56]   = Image[678];
    assign  image_0_635[55:48]   = Image[679];
    assign  image_0_635[47:40]   = Image[709];
    assign  image_0_635[39:32]   = Image[710];
    assign  image_0_635[31:24]   = Image[711];
    assign  image_0_635[23:16]   = Image[741];
    assign  image_0_635[15:8]    = Image[742];
    assign  image_0_635[7:0]     = Image[743];

    assign  image_0_636[71:64]   = Image[678];
    assign  image_0_636[63:56]   = Image[679];
    assign  image_0_636[55:48]   = Image[680];
    assign  image_0_636[47:40]   = Image[710];
    assign  image_0_636[39:32]   = Image[711];
    assign  image_0_636[31:24]   = Image[712];
    assign  image_0_636[23:16]   = Image[742];
    assign  image_0_636[15:8]    = Image[743];
    assign  image_0_636[7:0]     = Image[744];

    assign  image_0_637[71:64]   = Image[679];
    assign  image_0_637[63:56]   = Image[680];
    assign  image_0_637[55:48]   = Image[681];
    assign  image_0_637[47:40]   = Image[711];
    assign  image_0_637[39:32]   = Image[712];
    assign  image_0_637[31:24]   = Image[713];
    assign  image_0_637[23:16]   = Image[743];
    assign  image_0_637[15:8]    = Image[744];
    assign  image_0_637[7:0]     = Image[745];

    assign  image_0_638[71:64]   = Image[680];
    assign  image_0_638[63:56]   = Image[681];
    assign  image_0_638[55:48]   = Image[682];
    assign  image_0_638[47:40]   = Image[712];
    assign  image_0_638[39:32]   = Image[713];
    assign  image_0_638[31:24]   = Image[714];
    assign  image_0_638[23:16]   = Image[744];
    assign  image_0_638[15:8]    = Image[745];
    assign  image_0_638[7:0]     = Image[746];

    assign  image_0_639[71:64]   = Image[681];
    assign  image_0_639[63:56]   = Image[682];
    assign  image_0_639[55:48]   = Image[683];
    assign  image_0_639[47:40]   = Image[713];
    assign  image_0_639[39:32]   = Image[714];
    assign  image_0_639[31:24]   = Image[715];
    assign  image_0_639[23:16]   = Image[745];
    assign  image_0_639[15:8]    = Image[746];
    assign  image_0_639[7:0]     = Image[747];

    assign  image_0_640[71:64]   = Image[682];
    assign  image_0_640[63:56]   = Image[683];
    assign  image_0_640[55:48]   = Image[684];
    assign  image_0_640[47:40]   = Image[714];
    assign  image_0_640[39:32]   = Image[715];
    assign  image_0_640[31:24]   = Image[716];
    assign  image_0_640[23:16]   = Image[746];
    assign  image_0_640[15:8]    = Image[747];
    assign  image_0_640[7:0]     = Image[748];

    assign  image_0_641[71:64]   = Image[683];
    assign  image_0_641[63:56]   = Image[684];
    assign  image_0_641[55:48]   = Image[685];
    assign  image_0_641[47:40]   = Image[715];
    assign  image_0_641[39:32]   = Image[716];
    assign  image_0_641[31:24]   = Image[717];
    assign  image_0_641[23:16]   = Image[747];
    assign  image_0_641[15:8]    = Image[748];
    assign  image_0_641[7:0]     = Image[749];

    assign  image_0_642[71:64]   = Image[684];
    assign  image_0_642[63:56]   = Image[685];
    assign  image_0_642[55:48]   = Image[686];
    assign  image_0_642[47:40]   = Image[716];
    assign  image_0_642[39:32]   = Image[717];
    assign  image_0_642[31:24]   = Image[718];
    assign  image_0_642[23:16]   = Image[748];
    assign  image_0_642[15:8]    = Image[749];
    assign  image_0_642[7:0]     = Image[750];

    assign  image_0_643[71:64]   = Image[685];
    assign  image_0_643[63:56]   = Image[686];
    assign  image_0_643[55:48]   = Image[687];
    assign  image_0_643[47:40]   = Image[717];
    assign  image_0_643[39:32]   = Image[718];
    assign  image_0_643[31:24]   = Image[719];
    assign  image_0_643[23:16]   = Image[749];
    assign  image_0_643[15:8]    = Image[750];
    assign  image_0_643[7:0]     = Image[751];

    assign  image_0_644[71:64]   = Image[686];
    assign  image_0_644[63:56]   = Image[687];
    assign  image_0_644[55:48]   = Image[688];
    assign  image_0_644[47:40]   = Image[718];
    assign  image_0_644[39:32]   = Image[719];
    assign  image_0_644[31:24]   = Image[720];
    assign  image_0_644[23:16]   = Image[750];
    assign  image_0_644[15:8]    = Image[751];
    assign  image_0_644[7:0]     = Image[752];

    assign  image_0_645[71:64]   = Image[687];
    assign  image_0_645[63:56]   = Image[688];
    assign  image_0_645[55:48]   = Image[689];
    assign  image_0_645[47:40]   = Image[719];
    assign  image_0_645[39:32]   = Image[720];
    assign  image_0_645[31:24]   = Image[721];
    assign  image_0_645[23:16]   = Image[751];
    assign  image_0_645[15:8]    = Image[752];
    assign  image_0_645[7:0]     = Image[753];

    assign  image_0_646[71:64]   = Image[688];
    assign  image_0_646[63:56]   = Image[689];
    assign  image_0_646[55:48]   = Image[690];
    assign  image_0_646[47:40]   = Image[720];
    assign  image_0_646[39:32]   = Image[721];
    assign  image_0_646[31:24]   = Image[722];
    assign  image_0_646[23:16]   = Image[752];
    assign  image_0_646[15:8]    = Image[753];
    assign  image_0_646[7:0]     = Image[754];

    assign  image_0_647[71:64]   = Image[689];
    assign  image_0_647[63:56]   = Image[690];
    assign  image_0_647[55:48]   = Image[691];
    assign  image_0_647[47:40]   = Image[721];
    assign  image_0_647[39:32]   = Image[722];
    assign  image_0_647[31:24]   = Image[723];
    assign  image_0_647[23:16]   = Image[753];
    assign  image_0_647[15:8]    = Image[754];
    assign  image_0_647[7:0]     = Image[755];

    assign  image_0_648[71:64]   = Image[690];
    assign  image_0_648[63:56]   = Image[691];
    assign  image_0_648[55:48]   = Image[692];
    assign  image_0_648[47:40]   = Image[722];
    assign  image_0_648[39:32]   = Image[723];
    assign  image_0_648[31:24]   = Image[724];
    assign  image_0_648[23:16]   = Image[754];
    assign  image_0_648[15:8]    = Image[755];
    assign  image_0_648[7:0]     = Image[756];

    assign  image_0_649[71:64]   = Image[691];
    assign  image_0_649[63:56]   = Image[692];
    assign  image_0_649[55:48]   = Image[693];
    assign  image_0_649[47:40]   = Image[723];
    assign  image_0_649[39:32]   = Image[724];
    assign  image_0_649[31:24]   = Image[725];
    assign  image_0_649[23:16]   = Image[755];
    assign  image_0_649[15:8]    = Image[756];
    assign  image_0_649[7:0]     = Image[757];

    assign  image_0_650[71:64]   = Image[692];
    assign  image_0_650[63:56]   = Image[693];
    assign  image_0_650[55:48]   = Image[694];
    assign  image_0_650[47:40]   = Image[724];
    assign  image_0_650[39:32]   = Image[725];
    assign  image_0_650[31:24]   = Image[726];
    assign  image_0_650[23:16]   = Image[756];
    assign  image_0_650[15:8]    = Image[757];
    assign  image_0_650[7:0]     = Image[758];

    assign  image_0_651[71:64]   = Image[693];
    assign  image_0_651[63:56]   = Image[694];
    assign  image_0_651[55:48]   = Image[695];
    assign  image_0_651[47:40]   = Image[725];
    assign  image_0_651[39:32]   = Image[726];
    assign  image_0_651[31:24]   = Image[727];
    assign  image_0_651[23:16]   = Image[757];
    assign  image_0_651[15:8]    = Image[758];
    assign  image_0_651[7:0]     = Image[759];

    assign  image_0_652[71:64]   = Image[694];
    assign  image_0_652[63:56]   = Image[695];
    assign  image_0_652[55:48]   = Image[696];
    assign  image_0_652[47:40]   = Image[726];
    assign  image_0_652[39:32]   = Image[727];
    assign  image_0_652[31:24]   = Image[728];
    assign  image_0_652[23:16]   = Image[758];
    assign  image_0_652[15:8]    = Image[759];
    assign  image_0_652[7:0]     = Image[760];

    assign  image_0_653[71:64]   = Image[695];
    assign  image_0_653[63:56]   = Image[696];
    assign  image_0_653[55:48]   = Image[697];
    assign  image_0_653[47:40]   = Image[727];
    assign  image_0_653[39:32]   = Image[728];
    assign  image_0_653[31:24]   = Image[729];
    assign  image_0_653[23:16]   = Image[759];
    assign  image_0_653[15:8]    = Image[760];
    assign  image_0_653[7:0]     = Image[761];

    assign  image_0_654[71:64]   = Image[696];
    assign  image_0_654[63:56]   = Image[697];
    assign  image_0_654[55:48]   = Image[698];
    assign  image_0_654[47:40]   = Image[728];
    assign  image_0_654[39:32]   = Image[729];
    assign  image_0_654[31:24]   = Image[730];
    assign  image_0_654[23:16]   = Image[760];
    assign  image_0_654[15:8]    = Image[761];
    assign  image_0_654[7:0]     = Image[762];

    assign  image_0_655[71:64]   = Image[697];
    assign  image_0_655[63:56]   = Image[698];
    assign  image_0_655[55:48]   = Image[699];
    assign  image_0_655[47:40]   = Image[729];
    assign  image_0_655[39:32]   = Image[730];
    assign  image_0_655[31:24]   = Image[731];
    assign  image_0_655[23:16]   = Image[761];
    assign  image_0_655[15:8]    = Image[762];
    assign  image_0_655[7:0]     = Image[763];

    assign  image_0_656[71:64]   = Image[698];
    assign  image_0_656[63:56]   = Image[699];
    assign  image_0_656[55:48]   = Image[700];
    assign  image_0_656[47:40]   = Image[730];
    assign  image_0_656[39:32]   = Image[731];
    assign  image_0_656[31:24]   = Image[732];
    assign  image_0_656[23:16]   = Image[762];
    assign  image_0_656[15:8]    = Image[763];
    assign  image_0_656[7:0]     = Image[764];

    assign  image_0_657[71:64]   = Image[699];
    assign  image_0_657[63:56]   = Image[700];
    assign  image_0_657[55:48]   = Image[701];
    assign  image_0_657[47:40]   = Image[731];
    assign  image_0_657[39:32]   = Image[732];
    assign  image_0_657[31:24]   = Image[733];
    assign  image_0_657[23:16]   = Image[763];
    assign  image_0_657[15:8]    = Image[764];
    assign  image_0_657[7:0]     = Image[765];

    assign  image_0_658[71:64]   = Image[700];
    assign  image_0_658[63:56]   = Image[701];
    assign  image_0_658[55:48]   = Image[702];
    assign  image_0_658[47:40]   = Image[732];
    assign  image_0_658[39:32]   = Image[733];
    assign  image_0_658[31:24]   = Image[734];
    assign  image_0_658[23:16]   = Image[764];
    assign  image_0_658[15:8]    = Image[765];
    assign  image_0_658[7:0]     = Image[766];

    assign  image_0_659[71:64]   = Image[701];
    assign  image_0_659[63:56]   = Image[702];
    assign  image_0_659[55:48]   = Image[703];
    assign  image_0_659[47:40]   = Image[733];
    assign  image_0_659[39:32]   = Image[734];
    assign  image_0_659[31:24]   = Image[735];
    assign  image_0_659[23:16]   = Image[765];
    assign  image_0_659[15:8]    = Image[766];
    assign  image_0_659[7:0]     = Image[767];

    assign  image_0_660[71:64]   = Image[704];
    assign  image_0_660[63:56]   = Image[705];
    assign  image_0_660[55:48]   = Image[706];
    assign  image_0_660[47:40]   = Image[736];
    assign  image_0_660[39:32]   = Image[737];
    assign  image_0_660[31:24]   = Image[738];
    assign  image_0_660[23:16]   = Image[768];
    assign  image_0_660[15:8]    = Image[769];
    assign  image_0_660[7:0]     = Image[770];

    assign  image_0_661[71:64]   = Image[705];
    assign  image_0_661[63:56]   = Image[706];
    assign  image_0_661[55:48]   = Image[707];
    assign  image_0_661[47:40]   = Image[737];
    assign  image_0_661[39:32]   = Image[738];
    assign  image_0_661[31:24]   = Image[739];
    assign  image_0_661[23:16]   = Image[769];
    assign  image_0_661[15:8]    = Image[770];
    assign  image_0_661[7:0]     = Image[771];

    assign  image_0_662[71:64]   = Image[706];
    assign  image_0_662[63:56]   = Image[707];
    assign  image_0_662[55:48]   = Image[708];
    assign  image_0_662[47:40]   = Image[738];
    assign  image_0_662[39:32]   = Image[739];
    assign  image_0_662[31:24]   = Image[740];
    assign  image_0_662[23:16]   = Image[770];
    assign  image_0_662[15:8]    = Image[771];
    assign  image_0_662[7:0]     = Image[772];

    assign  image_0_663[71:64]   = Image[707];
    assign  image_0_663[63:56]   = Image[708];
    assign  image_0_663[55:48]   = Image[709];
    assign  image_0_663[47:40]   = Image[739];
    assign  image_0_663[39:32]   = Image[740];
    assign  image_0_663[31:24]   = Image[741];
    assign  image_0_663[23:16]   = Image[771];
    assign  image_0_663[15:8]    = Image[772];
    assign  image_0_663[7:0]     = Image[773];

    assign  image_0_664[71:64]   = Image[708];
    assign  image_0_664[63:56]   = Image[709];
    assign  image_0_664[55:48]   = Image[710];
    assign  image_0_664[47:40]   = Image[740];
    assign  image_0_664[39:32]   = Image[741];
    assign  image_0_664[31:24]   = Image[742];
    assign  image_0_664[23:16]   = Image[772];
    assign  image_0_664[15:8]    = Image[773];
    assign  image_0_664[7:0]     = Image[774];

    assign  image_0_665[71:64]   = Image[709];
    assign  image_0_665[63:56]   = Image[710];
    assign  image_0_665[55:48]   = Image[711];
    assign  image_0_665[47:40]   = Image[741];
    assign  image_0_665[39:32]   = Image[742];
    assign  image_0_665[31:24]   = Image[743];
    assign  image_0_665[23:16]   = Image[773];
    assign  image_0_665[15:8]    = Image[774];
    assign  image_0_665[7:0]     = Image[775];

    assign  image_0_666[71:64]   = Image[710];
    assign  image_0_666[63:56]   = Image[711];
    assign  image_0_666[55:48]   = Image[712];
    assign  image_0_666[47:40]   = Image[742];
    assign  image_0_666[39:32]   = Image[743];
    assign  image_0_666[31:24]   = Image[744];
    assign  image_0_666[23:16]   = Image[774];
    assign  image_0_666[15:8]    = Image[775];
    assign  image_0_666[7:0]     = Image[776];

    assign  image_0_667[71:64]   = Image[711];
    assign  image_0_667[63:56]   = Image[712];
    assign  image_0_667[55:48]   = Image[713];
    assign  image_0_667[47:40]   = Image[743];
    assign  image_0_667[39:32]   = Image[744];
    assign  image_0_667[31:24]   = Image[745];
    assign  image_0_667[23:16]   = Image[775];
    assign  image_0_667[15:8]    = Image[776];
    assign  image_0_667[7:0]     = Image[777];

    assign  image_0_668[71:64]   = Image[712];
    assign  image_0_668[63:56]   = Image[713];
    assign  image_0_668[55:48]   = Image[714];
    assign  image_0_668[47:40]   = Image[744];
    assign  image_0_668[39:32]   = Image[745];
    assign  image_0_668[31:24]   = Image[746];
    assign  image_0_668[23:16]   = Image[776];
    assign  image_0_668[15:8]    = Image[777];
    assign  image_0_668[7:0]     = Image[778];

    assign  image_0_669[71:64]   = Image[713];
    assign  image_0_669[63:56]   = Image[714];
    assign  image_0_669[55:48]   = Image[715];
    assign  image_0_669[47:40]   = Image[745];
    assign  image_0_669[39:32]   = Image[746];
    assign  image_0_669[31:24]   = Image[747];
    assign  image_0_669[23:16]   = Image[777];
    assign  image_0_669[15:8]    = Image[778];
    assign  image_0_669[7:0]     = Image[779];

    assign  image_0_670[71:64]   = Image[714];
    assign  image_0_670[63:56]   = Image[715];
    assign  image_0_670[55:48]   = Image[716];
    assign  image_0_670[47:40]   = Image[746];
    assign  image_0_670[39:32]   = Image[747];
    assign  image_0_670[31:24]   = Image[748];
    assign  image_0_670[23:16]   = Image[778];
    assign  image_0_670[15:8]    = Image[779];
    assign  image_0_670[7:0]     = Image[780];

    assign  image_0_671[71:64]   = Image[715];
    assign  image_0_671[63:56]   = Image[716];
    assign  image_0_671[55:48]   = Image[717];
    assign  image_0_671[47:40]   = Image[747];
    assign  image_0_671[39:32]   = Image[748];
    assign  image_0_671[31:24]   = Image[749];
    assign  image_0_671[23:16]   = Image[779];
    assign  image_0_671[15:8]    = Image[780];
    assign  image_0_671[7:0]     = Image[781];

    assign  image_0_672[71:64]   = Image[716];
    assign  image_0_672[63:56]   = Image[717];
    assign  image_0_672[55:48]   = Image[718];
    assign  image_0_672[47:40]   = Image[748];
    assign  image_0_672[39:32]   = Image[749];
    assign  image_0_672[31:24]   = Image[750];
    assign  image_0_672[23:16]   = Image[780];
    assign  image_0_672[15:8]    = Image[781];
    assign  image_0_672[7:0]     = Image[782];

    assign  image_0_673[71:64]   = Image[717];
    assign  image_0_673[63:56]   = Image[718];
    assign  image_0_673[55:48]   = Image[719];
    assign  image_0_673[47:40]   = Image[749];
    assign  image_0_673[39:32]   = Image[750];
    assign  image_0_673[31:24]   = Image[751];
    assign  image_0_673[23:16]   = Image[781];
    assign  image_0_673[15:8]    = Image[782];
    assign  image_0_673[7:0]     = Image[783];

    assign  image_0_674[71:64]   = Image[718];
    assign  image_0_674[63:56]   = Image[719];
    assign  image_0_674[55:48]   = Image[720];
    assign  image_0_674[47:40]   = Image[750];
    assign  image_0_674[39:32]   = Image[751];
    assign  image_0_674[31:24]   = Image[752];
    assign  image_0_674[23:16]   = Image[782];
    assign  image_0_674[15:8]    = Image[783];
    assign  image_0_674[7:0]     = Image[784];

    assign  image_0_675[71:64]   = Image[719];
    assign  image_0_675[63:56]   = Image[720];
    assign  image_0_675[55:48]   = Image[721];
    assign  image_0_675[47:40]   = Image[751];
    assign  image_0_675[39:32]   = Image[752];
    assign  image_0_675[31:24]   = Image[753];
    assign  image_0_675[23:16]   = Image[783];
    assign  image_0_675[15:8]    = Image[784];
    assign  image_0_675[7:0]     = Image[785];

    assign  image_0_676[71:64]   = Image[720];
    assign  image_0_676[63:56]   = Image[721];
    assign  image_0_676[55:48]   = Image[722];
    assign  image_0_676[47:40]   = Image[752];
    assign  image_0_676[39:32]   = Image[753];
    assign  image_0_676[31:24]   = Image[754];
    assign  image_0_676[23:16]   = Image[784];
    assign  image_0_676[15:8]    = Image[785];
    assign  image_0_676[7:0]     = Image[786];

    assign  image_0_677[71:64]   = Image[721];
    assign  image_0_677[63:56]   = Image[722];
    assign  image_0_677[55:48]   = Image[723];
    assign  image_0_677[47:40]   = Image[753];
    assign  image_0_677[39:32]   = Image[754];
    assign  image_0_677[31:24]   = Image[755];
    assign  image_0_677[23:16]   = Image[785];
    assign  image_0_677[15:8]    = Image[786];
    assign  image_0_677[7:0]     = Image[787];

    assign  image_0_678[71:64]   = Image[722];
    assign  image_0_678[63:56]   = Image[723];
    assign  image_0_678[55:48]   = Image[724];
    assign  image_0_678[47:40]   = Image[754];
    assign  image_0_678[39:32]   = Image[755];
    assign  image_0_678[31:24]   = Image[756];
    assign  image_0_678[23:16]   = Image[786];
    assign  image_0_678[15:8]    = Image[787];
    assign  image_0_678[7:0]     = Image[788];

    assign  image_0_679[71:64]   = Image[723];
    assign  image_0_679[63:56]   = Image[724];
    assign  image_0_679[55:48]   = Image[725];
    assign  image_0_679[47:40]   = Image[755];
    assign  image_0_679[39:32]   = Image[756];
    assign  image_0_679[31:24]   = Image[757];
    assign  image_0_679[23:16]   = Image[787];
    assign  image_0_679[15:8]    = Image[788];
    assign  image_0_679[7:0]     = Image[789];

    assign  image_0_680[71:64]   = Image[724];
    assign  image_0_680[63:56]   = Image[725];
    assign  image_0_680[55:48]   = Image[726];
    assign  image_0_680[47:40]   = Image[756];
    assign  image_0_680[39:32]   = Image[757];
    assign  image_0_680[31:24]   = Image[758];
    assign  image_0_680[23:16]   = Image[788];
    assign  image_0_680[15:8]    = Image[789];
    assign  image_0_680[7:0]     = Image[790];

    assign  image_0_681[71:64]   = Image[725];
    assign  image_0_681[63:56]   = Image[726];
    assign  image_0_681[55:48]   = Image[727];
    assign  image_0_681[47:40]   = Image[757];
    assign  image_0_681[39:32]   = Image[758];
    assign  image_0_681[31:24]   = Image[759];
    assign  image_0_681[23:16]   = Image[789];
    assign  image_0_681[15:8]    = Image[790];
    assign  image_0_681[7:0]     = Image[791];

    assign  image_0_682[71:64]   = Image[726];
    assign  image_0_682[63:56]   = Image[727];
    assign  image_0_682[55:48]   = Image[728];
    assign  image_0_682[47:40]   = Image[758];
    assign  image_0_682[39:32]   = Image[759];
    assign  image_0_682[31:24]   = Image[760];
    assign  image_0_682[23:16]   = Image[790];
    assign  image_0_682[15:8]    = Image[791];
    assign  image_0_682[7:0]     = Image[792];

    assign  image_0_683[71:64]   = Image[727];
    assign  image_0_683[63:56]   = Image[728];
    assign  image_0_683[55:48]   = Image[729];
    assign  image_0_683[47:40]   = Image[759];
    assign  image_0_683[39:32]   = Image[760];
    assign  image_0_683[31:24]   = Image[761];
    assign  image_0_683[23:16]   = Image[791];
    assign  image_0_683[15:8]    = Image[792];
    assign  image_0_683[7:0]     = Image[793];

    assign  image_0_684[71:64]   = Image[728];
    assign  image_0_684[63:56]   = Image[729];
    assign  image_0_684[55:48]   = Image[730];
    assign  image_0_684[47:40]   = Image[760];
    assign  image_0_684[39:32]   = Image[761];
    assign  image_0_684[31:24]   = Image[762];
    assign  image_0_684[23:16]   = Image[792];
    assign  image_0_684[15:8]    = Image[793];
    assign  image_0_684[7:0]     = Image[794];

    assign  image_0_685[71:64]   = Image[729];
    assign  image_0_685[63:56]   = Image[730];
    assign  image_0_685[55:48]   = Image[731];
    assign  image_0_685[47:40]   = Image[761];
    assign  image_0_685[39:32]   = Image[762];
    assign  image_0_685[31:24]   = Image[763];
    assign  image_0_685[23:16]   = Image[793];
    assign  image_0_685[15:8]    = Image[794];
    assign  image_0_685[7:0]     = Image[795];

    assign  image_0_686[71:64]   = Image[730];
    assign  image_0_686[63:56]   = Image[731];
    assign  image_0_686[55:48]   = Image[732];
    assign  image_0_686[47:40]   = Image[762];
    assign  image_0_686[39:32]   = Image[763];
    assign  image_0_686[31:24]   = Image[764];
    assign  image_0_686[23:16]   = Image[794];
    assign  image_0_686[15:8]    = Image[795];
    assign  image_0_686[7:0]     = Image[796];

    assign  image_0_687[71:64]   = Image[731];
    assign  image_0_687[63:56]   = Image[732];
    assign  image_0_687[55:48]   = Image[733];
    assign  image_0_687[47:40]   = Image[763];
    assign  image_0_687[39:32]   = Image[764];
    assign  image_0_687[31:24]   = Image[765];
    assign  image_0_687[23:16]   = Image[795];
    assign  image_0_687[15:8]    = Image[796];
    assign  image_0_687[7:0]     = Image[797];

    assign  image_0_688[71:64]   = Image[732];
    assign  image_0_688[63:56]   = Image[733];
    assign  image_0_688[55:48]   = Image[734];
    assign  image_0_688[47:40]   = Image[764];
    assign  image_0_688[39:32]   = Image[765];
    assign  image_0_688[31:24]   = Image[766];
    assign  image_0_688[23:16]   = Image[796];
    assign  image_0_688[15:8]    = Image[797];
    assign  image_0_688[7:0]     = Image[798];

    assign  image_0_689[71:64]   = Image[733];
    assign  image_0_689[63:56]   = Image[734];
    assign  image_0_689[55:48]   = Image[735];
    assign  image_0_689[47:40]   = Image[765];
    assign  image_0_689[39:32]   = Image[766];
    assign  image_0_689[31:24]   = Image[767];
    assign  image_0_689[23:16]   = Image[797];
    assign  image_0_689[15:8]    = Image[798];
    assign  image_0_689[7:0]     = Image[799];

    assign  image_0_690[71:64]   = Image[736];
    assign  image_0_690[63:56]   = Image[737];
    assign  image_0_690[55:48]   = Image[738];
    assign  image_0_690[47:40]   = Image[768];
    assign  image_0_690[39:32]   = Image[769];
    assign  image_0_690[31:24]   = Image[770];
    assign  image_0_690[23:16]   = Image[800];
    assign  image_0_690[15:8]    = Image[801];
    assign  image_0_690[7:0]     = Image[802];

    assign  image_0_691[71:64]   = Image[737];
    assign  image_0_691[63:56]   = Image[738];
    assign  image_0_691[55:48]   = Image[739];
    assign  image_0_691[47:40]   = Image[769];
    assign  image_0_691[39:32]   = Image[770];
    assign  image_0_691[31:24]   = Image[771];
    assign  image_0_691[23:16]   = Image[801];
    assign  image_0_691[15:8]    = Image[802];
    assign  image_0_691[7:0]     = Image[803];

    assign  image_0_692[71:64]   = Image[738];
    assign  image_0_692[63:56]   = Image[739];
    assign  image_0_692[55:48]   = Image[740];
    assign  image_0_692[47:40]   = Image[770];
    assign  image_0_692[39:32]   = Image[771];
    assign  image_0_692[31:24]   = Image[772];
    assign  image_0_692[23:16]   = Image[802];
    assign  image_0_692[15:8]    = Image[803];
    assign  image_0_692[7:0]     = Image[804];

    assign  image_0_693[71:64]   = Image[739];
    assign  image_0_693[63:56]   = Image[740];
    assign  image_0_693[55:48]   = Image[741];
    assign  image_0_693[47:40]   = Image[771];
    assign  image_0_693[39:32]   = Image[772];
    assign  image_0_693[31:24]   = Image[773];
    assign  image_0_693[23:16]   = Image[803];
    assign  image_0_693[15:8]    = Image[804];
    assign  image_0_693[7:0]     = Image[805];

    assign  image_0_694[71:64]   = Image[740];
    assign  image_0_694[63:56]   = Image[741];
    assign  image_0_694[55:48]   = Image[742];
    assign  image_0_694[47:40]   = Image[772];
    assign  image_0_694[39:32]   = Image[773];
    assign  image_0_694[31:24]   = Image[774];
    assign  image_0_694[23:16]   = Image[804];
    assign  image_0_694[15:8]    = Image[805];
    assign  image_0_694[7:0]     = Image[806];

    assign  image_0_695[71:64]   = Image[741];
    assign  image_0_695[63:56]   = Image[742];
    assign  image_0_695[55:48]   = Image[743];
    assign  image_0_695[47:40]   = Image[773];
    assign  image_0_695[39:32]   = Image[774];
    assign  image_0_695[31:24]   = Image[775];
    assign  image_0_695[23:16]   = Image[805];
    assign  image_0_695[15:8]    = Image[806];
    assign  image_0_695[7:0]     = Image[807];

    assign  image_0_696[71:64]   = Image[742];
    assign  image_0_696[63:56]   = Image[743];
    assign  image_0_696[55:48]   = Image[744];
    assign  image_0_696[47:40]   = Image[774];
    assign  image_0_696[39:32]   = Image[775];
    assign  image_0_696[31:24]   = Image[776];
    assign  image_0_696[23:16]   = Image[806];
    assign  image_0_696[15:8]    = Image[807];
    assign  image_0_696[7:0]     = Image[808];

    assign  image_0_697[71:64]   = Image[743];
    assign  image_0_697[63:56]   = Image[744];
    assign  image_0_697[55:48]   = Image[745];
    assign  image_0_697[47:40]   = Image[775];
    assign  image_0_697[39:32]   = Image[776];
    assign  image_0_697[31:24]   = Image[777];
    assign  image_0_697[23:16]   = Image[807];
    assign  image_0_697[15:8]    = Image[808];
    assign  image_0_697[7:0]     = Image[809];

    assign  image_0_698[71:64]   = Image[744];
    assign  image_0_698[63:56]   = Image[745];
    assign  image_0_698[55:48]   = Image[746];
    assign  image_0_698[47:40]   = Image[776];
    assign  image_0_698[39:32]   = Image[777];
    assign  image_0_698[31:24]   = Image[778];
    assign  image_0_698[23:16]   = Image[808];
    assign  image_0_698[15:8]    = Image[809];
    assign  image_0_698[7:0]     = Image[810];

    assign  image_0_699[71:64]   = Image[745];
    assign  image_0_699[63:56]   = Image[746];
    assign  image_0_699[55:48]   = Image[747];
    assign  image_0_699[47:40]   = Image[777];
    assign  image_0_699[39:32]   = Image[778];
    assign  image_0_699[31:24]   = Image[779];
    assign  image_0_699[23:16]   = Image[809];
    assign  image_0_699[15:8]    = Image[810];
    assign  image_0_699[7:0]     = Image[811];

    assign  image_0_700[71:64]   = Image[746];
    assign  image_0_700[63:56]   = Image[747];
    assign  image_0_700[55:48]   = Image[748];
    assign  image_0_700[47:40]   = Image[778];
    assign  image_0_700[39:32]   = Image[779];
    assign  image_0_700[31:24]   = Image[780];
    assign  image_0_700[23:16]   = Image[810];
    assign  image_0_700[15:8]    = Image[811];
    assign  image_0_700[7:0]     = Image[812];

    assign  image_0_701[71:64]   = Image[747];
    assign  image_0_701[63:56]   = Image[748];
    assign  image_0_701[55:48]   = Image[749];
    assign  image_0_701[47:40]   = Image[779];
    assign  image_0_701[39:32]   = Image[780];
    assign  image_0_701[31:24]   = Image[781];
    assign  image_0_701[23:16]   = Image[811];
    assign  image_0_701[15:8]    = Image[812];
    assign  image_0_701[7:0]     = Image[813];

    assign  image_0_702[71:64]   = Image[748];
    assign  image_0_702[63:56]   = Image[749];
    assign  image_0_702[55:48]   = Image[750];
    assign  image_0_702[47:40]   = Image[780];
    assign  image_0_702[39:32]   = Image[781];
    assign  image_0_702[31:24]   = Image[782];
    assign  image_0_702[23:16]   = Image[812];
    assign  image_0_702[15:8]    = Image[813];
    assign  image_0_702[7:0]     = Image[814];

    assign  image_0_703[71:64]   = Image[749];
    assign  image_0_703[63:56]   = Image[750];
    assign  image_0_703[55:48]   = Image[751];
    assign  image_0_703[47:40]   = Image[781];
    assign  image_0_703[39:32]   = Image[782];
    assign  image_0_703[31:24]   = Image[783];
    assign  image_0_703[23:16]   = Image[813];
    assign  image_0_703[15:8]    = Image[814];
    assign  image_0_703[7:0]     = Image[815];

    assign  image_0_704[71:64]   = Image[750];
    assign  image_0_704[63:56]   = Image[751];
    assign  image_0_704[55:48]   = Image[752];
    assign  image_0_704[47:40]   = Image[782];
    assign  image_0_704[39:32]   = Image[783];
    assign  image_0_704[31:24]   = Image[784];
    assign  image_0_704[23:16]   = Image[814];
    assign  image_0_704[15:8]    = Image[815];
    assign  image_0_704[7:0]     = Image[816];

    assign  image_0_705[71:64]   = Image[751];
    assign  image_0_705[63:56]   = Image[752];
    assign  image_0_705[55:48]   = Image[753];
    assign  image_0_705[47:40]   = Image[783];
    assign  image_0_705[39:32]   = Image[784];
    assign  image_0_705[31:24]   = Image[785];
    assign  image_0_705[23:16]   = Image[815];
    assign  image_0_705[15:8]    = Image[816];
    assign  image_0_705[7:0]     = Image[817];

    assign  image_0_706[71:64]   = Image[752];
    assign  image_0_706[63:56]   = Image[753];
    assign  image_0_706[55:48]   = Image[754];
    assign  image_0_706[47:40]   = Image[784];
    assign  image_0_706[39:32]   = Image[785];
    assign  image_0_706[31:24]   = Image[786];
    assign  image_0_706[23:16]   = Image[816];
    assign  image_0_706[15:8]    = Image[817];
    assign  image_0_706[7:0]     = Image[818];

    assign  image_0_707[71:64]   = Image[753];
    assign  image_0_707[63:56]   = Image[754];
    assign  image_0_707[55:48]   = Image[755];
    assign  image_0_707[47:40]   = Image[785];
    assign  image_0_707[39:32]   = Image[786];
    assign  image_0_707[31:24]   = Image[787];
    assign  image_0_707[23:16]   = Image[817];
    assign  image_0_707[15:8]    = Image[818];
    assign  image_0_707[7:0]     = Image[819];

    assign  image_0_708[71:64]   = Image[754];
    assign  image_0_708[63:56]   = Image[755];
    assign  image_0_708[55:48]   = Image[756];
    assign  image_0_708[47:40]   = Image[786];
    assign  image_0_708[39:32]   = Image[787];
    assign  image_0_708[31:24]   = Image[788];
    assign  image_0_708[23:16]   = Image[818];
    assign  image_0_708[15:8]    = Image[819];
    assign  image_0_708[7:0]     = Image[820];

    assign  image_0_709[71:64]   = Image[755];
    assign  image_0_709[63:56]   = Image[756];
    assign  image_0_709[55:48]   = Image[757];
    assign  image_0_709[47:40]   = Image[787];
    assign  image_0_709[39:32]   = Image[788];
    assign  image_0_709[31:24]   = Image[789];
    assign  image_0_709[23:16]   = Image[819];
    assign  image_0_709[15:8]    = Image[820];
    assign  image_0_709[7:0]     = Image[821];

    assign  image_0_710[71:64]   = Image[756];
    assign  image_0_710[63:56]   = Image[757];
    assign  image_0_710[55:48]   = Image[758];
    assign  image_0_710[47:40]   = Image[788];
    assign  image_0_710[39:32]   = Image[789];
    assign  image_0_710[31:24]   = Image[790];
    assign  image_0_710[23:16]   = Image[820];
    assign  image_0_710[15:8]    = Image[821];
    assign  image_0_710[7:0]     = Image[822];

    assign  image_0_711[71:64]   = Image[757];
    assign  image_0_711[63:56]   = Image[758];
    assign  image_0_711[55:48]   = Image[759];
    assign  image_0_711[47:40]   = Image[789];
    assign  image_0_711[39:32]   = Image[790];
    assign  image_0_711[31:24]   = Image[791];
    assign  image_0_711[23:16]   = Image[821];
    assign  image_0_711[15:8]    = Image[822];
    assign  image_0_711[7:0]     = Image[823];

    assign  image_0_712[71:64]   = Image[758];
    assign  image_0_712[63:56]   = Image[759];
    assign  image_0_712[55:48]   = Image[760];
    assign  image_0_712[47:40]   = Image[790];
    assign  image_0_712[39:32]   = Image[791];
    assign  image_0_712[31:24]   = Image[792];
    assign  image_0_712[23:16]   = Image[822];
    assign  image_0_712[15:8]    = Image[823];
    assign  image_0_712[7:0]     = Image[824];

    assign  image_0_713[71:64]   = Image[759];
    assign  image_0_713[63:56]   = Image[760];
    assign  image_0_713[55:48]   = Image[761];
    assign  image_0_713[47:40]   = Image[791];
    assign  image_0_713[39:32]   = Image[792];
    assign  image_0_713[31:24]   = Image[793];
    assign  image_0_713[23:16]   = Image[823];
    assign  image_0_713[15:8]    = Image[824];
    assign  image_0_713[7:0]     = Image[825];

    assign  image_0_714[71:64]   = Image[760];
    assign  image_0_714[63:56]   = Image[761];
    assign  image_0_714[55:48]   = Image[762];
    assign  image_0_714[47:40]   = Image[792];
    assign  image_0_714[39:32]   = Image[793];
    assign  image_0_714[31:24]   = Image[794];
    assign  image_0_714[23:16]   = Image[824];
    assign  image_0_714[15:8]    = Image[825];
    assign  image_0_714[7:0]     = Image[826];

    assign  image_0_715[71:64]   = Image[761];
    assign  image_0_715[63:56]   = Image[762];
    assign  image_0_715[55:48]   = Image[763];
    assign  image_0_715[47:40]   = Image[793];
    assign  image_0_715[39:32]   = Image[794];
    assign  image_0_715[31:24]   = Image[795];
    assign  image_0_715[23:16]   = Image[825];
    assign  image_0_715[15:8]    = Image[826];
    assign  image_0_715[7:0]     = Image[827];

    assign  image_0_716[71:64]   = Image[762];
    assign  image_0_716[63:56]   = Image[763];
    assign  image_0_716[55:48]   = Image[764];
    assign  image_0_716[47:40]   = Image[794];
    assign  image_0_716[39:32]   = Image[795];
    assign  image_0_716[31:24]   = Image[796];
    assign  image_0_716[23:16]   = Image[826];
    assign  image_0_716[15:8]    = Image[827];
    assign  image_0_716[7:0]     = Image[828];

    assign  image_0_717[71:64]   = Image[763];
    assign  image_0_717[63:56]   = Image[764];
    assign  image_0_717[55:48]   = Image[765];
    assign  image_0_717[47:40]   = Image[795];
    assign  image_0_717[39:32]   = Image[796];
    assign  image_0_717[31:24]   = Image[797];
    assign  image_0_717[23:16]   = Image[827];
    assign  image_0_717[15:8]    = Image[828];
    assign  image_0_717[7:0]     = Image[829];

    assign  image_0_718[71:64]   = Image[764];
    assign  image_0_718[63:56]   = Image[765];
    assign  image_0_718[55:48]   = Image[766];
    assign  image_0_718[47:40]   = Image[796];
    assign  image_0_718[39:32]   = Image[797];
    assign  image_0_718[31:24]   = Image[798];
    assign  image_0_718[23:16]   = Image[828];
    assign  image_0_718[15:8]    = Image[829];
    assign  image_0_718[7:0]     = Image[830];

    assign  image_0_719[71:64]   = Image[765];
    assign  image_0_719[63:56]   = Image[766];
    assign  image_0_719[55:48]   = Image[767];
    assign  image_0_719[47:40]   = Image[797];
    assign  image_0_719[39:32]   = Image[798];
    assign  image_0_719[31:24]   = Image[799];
    assign  image_0_719[23:16]   = Image[829];
    assign  image_0_719[15:8]    = Image[830];
    assign  image_0_719[7:0]     = Image[831];

    assign  image_0_720[71:64]   = Image[768];
    assign  image_0_720[63:56]   = Image[769];
    assign  image_0_720[55:48]   = Image[770];
    assign  image_0_720[47:40]   = Image[800];
    assign  image_0_720[39:32]   = Image[801];
    assign  image_0_720[31:24]   = Image[802];
    assign  image_0_720[23:16]   = Image[832];
    assign  image_0_720[15:8]    = Image[833];
    assign  image_0_720[7:0]     = Image[834];

    assign  image_0_721[71:64]   = Image[769];
    assign  image_0_721[63:56]   = Image[770];
    assign  image_0_721[55:48]   = Image[771];
    assign  image_0_721[47:40]   = Image[801];
    assign  image_0_721[39:32]   = Image[802];
    assign  image_0_721[31:24]   = Image[803];
    assign  image_0_721[23:16]   = Image[833];
    assign  image_0_721[15:8]    = Image[834];
    assign  image_0_721[7:0]     = Image[835];

    assign  image_0_722[71:64]   = Image[770];
    assign  image_0_722[63:56]   = Image[771];
    assign  image_0_722[55:48]   = Image[772];
    assign  image_0_722[47:40]   = Image[802];
    assign  image_0_722[39:32]   = Image[803];
    assign  image_0_722[31:24]   = Image[804];
    assign  image_0_722[23:16]   = Image[834];
    assign  image_0_722[15:8]    = Image[835];
    assign  image_0_722[7:0]     = Image[836];

    assign  image_0_723[71:64]   = Image[771];
    assign  image_0_723[63:56]   = Image[772];
    assign  image_0_723[55:48]   = Image[773];
    assign  image_0_723[47:40]   = Image[803];
    assign  image_0_723[39:32]   = Image[804];
    assign  image_0_723[31:24]   = Image[805];
    assign  image_0_723[23:16]   = Image[835];
    assign  image_0_723[15:8]    = Image[836];
    assign  image_0_723[7:0]     = Image[837];

    assign  image_0_724[71:64]   = Image[772];
    assign  image_0_724[63:56]   = Image[773];
    assign  image_0_724[55:48]   = Image[774];
    assign  image_0_724[47:40]   = Image[804];
    assign  image_0_724[39:32]   = Image[805];
    assign  image_0_724[31:24]   = Image[806];
    assign  image_0_724[23:16]   = Image[836];
    assign  image_0_724[15:8]    = Image[837];
    assign  image_0_724[7:0]     = Image[838];

    assign  image_0_725[71:64]   = Image[773];
    assign  image_0_725[63:56]   = Image[774];
    assign  image_0_725[55:48]   = Image[775];
    assign  image_0_725[47:40]   = Image[805];
    assign  image_0_725[39:32]   = Image[806];
    assign  image_0_725[31:24]   = Image[807];
    assign  image_0_725[23:16]   = Image[837];
    assign  image_0_725[15:8]    = Image[838];
    assign  image_0_725[7:0]     = Image[839];

    assign  image_0_726[71:64]   = Image[774];
    assign  image_0_726[63:56]   = Image[775];
    assign  image_0_726[55:48]   = Image[776];
    assign  image_0_726[47:40]   = Image[806];
    assign  image_0_726[39:32]   = Image[807];
    assign  image_0_726[31:24]   = Image[808];
    assign  image_0_726[23:16]   = Image[838];
    assign  image_0_726[15:8]    = Image[839];
    assign  image_0_726[7:0]     = Image[840];

    assign  image_0_727[71:64]   = Image[775];
    assign  image_0_727[63:56]   = Image[776];
    assign  image_0_727[55:48]   = Image[777];
    assign  image_0_727[47:40]   = Image[807];
    assign  image_0_727[39:32]   = Image[808];
    assign  image_0_727[31:24]   = Image[809];
    assign  image_0_727[23:16]   = Image[839];
    assign  image_0_727[15:8]    = Image[840];
    assign  image_0_727[7:0]     = Image[841];

    assign  image_0_728[71:64]   = Image[776];
    assign  image_0_728[63:56]   = Image[777];
    assign  image_0_728[55:48]   = Image[778];
    assign  image_0_728[47:40]   = Image[808];
    assign  image_0_728[39:32]   = Image[809];
    assign  image_0_728[31:24]   = Image[810];
    assign  image_0_728[23:16]   = Image[840];
    assign  image_0_728[15:8]    = Image[841];
    assign  image_0_728[7:0]     = Image[842];

    assign  image_0_729[71:64]   = Image[777];
    assign  image_0_729[63:56]   = Image[778];
    assign  image_0_729[55:48]   = Image[779];
    assign  image_0_729[47:40]   = Image[809];
    assign  image_0_729[39:32]   = Image[810];
    assign  image_0_729[31:24]   = Image[811];
    assign  image_0_729[23:16]   = Image[841];
    assign  image_0_729[15:8]    = Image[842];
    assign  image_0_729[7:0]     = Image[843];

    assign  image_0_730[71:64]   = Image[778];
    assign  image_0_730[63:56]   = Image[779];
    assign  image_0_730[55:48]   = Image[780];
    assign  image_0_730[47:40]   = Image[810];
    assign  image_0_730[39:32]   = Image[811];
    assign  image_0_730[31:24]   = Image[812];
    assign  image_0_730[23:16]   = Image[842];
    assign  image_0_730[15:8]    = Image[843];
    assign  image_0_730[7:0]     = Image[844];

    assign  image_0_731[71:64]   = Image[779];
    assign  image_0_731[63:56]   = Image[780];
    assign  image_0_731[55:48]   = Image[781];
    assign  image_0_731[47:40]   = Image[811];
    assign  image_0_731[39:32]   = Image[812];
    assign  image_0_731[31:24]   = Image[813];
    assign  image_0_731[23:16]   = Image[843];
    assign  image_0_731[15:8]    = Image[844];
    assign  image_0_731[7:0]     = Image[845];

    assign  image_0_732[71:64]   = Image[780];
    assign  image_0_732[63:56]   = Image[781];
    assign  image_0_732[55:48]   = Image[782];
    assign  image_0_732[47:40]   = Image[812];
    assign  image_0_732[39:32]   = Image[813];
    assign  image_0_732[31:24]   = Image[814];
    assign  image_0_732[23:16]   = Image[844];
    assign  image_0_732[15:8]    = Image[845];
    assign  image_0_732[7:0]     = Image[846];

    assign  image_0_733[71:64]   = Image[781];
    assign  image_0_733[63:56]   = Image[782];
    assign  image_0_733[55:48]   = Image[783];
    assign  image_0_733[47:40]   = Image[813];
    assign  image_0_733[39:32]   = Image[814];
    assign  image_0_733[31:24]   = Image[815];
    assign  image_0_733[23:16]   = Image[845];
    assign  image_0_733[15:8]    = Image[846];
    assign  image_0_733[7:0]     = Image[847];

    assign  image_0_734[71:64]   = Image[782];
    assign  image_0_734[63:56]   = Image[783];
    assign  image_0_734[55:48]   = Image[784];
    assign  image_0_734[47:40]   = Image[814];
    assign  image_0_734[39:32]   = Image[815];
    assign  image_0_734[31:24]   = Image[816];
    assign  image_0_734[23:16]   = Image[846];
    assign  image_0_734[15:8]    = Image[847];
    assign  image_0_734[7:0]     = Image[848];

    assign  image_0_735[71:64]   = Image[783];
    assign  image_0_735[63:56]   = Image[784];
    assign  image_0_735[55:48]   = Image[785];
    assign  image_0_735[47:40]   = Image[815];
    assign  image_0_735[39:32]   = Image[816];
    assign  image_0_735[31:24]   = Image[817];
    assign  image_0_735[23:16]   = Image[847];
    assign  image_0_735[15:8]    = Image[848];
    assign  image_0_735[7:0]     = Image[849];

    assign  image_0_736[71:64]   = Image[784];
    assign  image_0_736[63:56]   = Image[785];
    assign  image_0_736[55:48]   = Image[786];
    assign  image_0_736[47:40]   = Image[816];
    assign  image_0_736[39:32]   = Image[817];
    assign  image_0_736[31:24]   = Image[818];
    assign  image_0_736[23:16]   = Image[848];
    assign  image_0_736[15:8]    = Image[849];
    assign  image_0_736[7:0]     = Image[850];

    assign  image_0_737[71:64]   = Image[785];
    assign  image_0_737[63:56]   = Image[786];
    assign  image_0_737[55:48]   = Image[787];
    assign  image_0_737[47:40]   = Image[817];
    assign  image_0_737[39:32]   = Image[818];
    assign  image_0_737[31:24]   = Image[819];
    assign  image_0_737[23:16]   = Image[849];
    assign  image_0_737[15:8]    = Image[850];
    assign  image_0_737[7:0]     = Image[851];

    assign  image_0_738[71:64]   = Image[786];
    assign  image_0_738[63:56]   = Image[787];
    assign  image_0_738[55:48]   = Image[788];
    assign  image_0_738[47:40]   = Image[818];
    assign  image_0_738[39:32]   = Image[819];
    assign  image_0_738[31:24]   = Image[820];
    assign  image_0_738[23:16]   = Image[850];
    assign  image_0_738[15:8]    = Image[851];
    assign  image_0_738[7:0]     = Image[852];

    assign  image_0_739[71:64]   = Image[787];
    assign  image_0_739[63:56]   = Image[788];
    assign  image_0_739[55:48]   = Image[789];
    assign  image_0_739[47:40]   = Image[819];
    assign  image_0_739[39:32]   = Image[820];
    assign  image_0_739[31:24]   = Image[821];
    assign  image_0_739[23:16]   = Image[851];
    assign  image_0_739[15:8]    = Image[852];
    assign  image_0_739[7:0]     = Image[853];

    assign  image_0_740[71:64]   = Image[788];
    assign  image_0_740[63:56]   = Image[789];
    assign  image_0_740[55:48]   = Image[790];
    assign  image_0_740[47:40]   = Image[820];
    assign  image_0_740[39:32]   = Image[821];
    assign  image_0_740[31:24]   = Image[822];
    assign  image_0_740[23:16]   = Image[852];
    assign  image_0_740[15:8]    = Image[853];
    assign  image_0_740[7:0]     = Image[854];

    assign  image_0_741[71:64]   = Image[789];
    assign  image_0_741[63:56]   = Image[790];
    assign  image_0_741[55:48]   = Image[791];
    assign  image_0_741[47:40]   = Image[821];
    assign  image_0_741[39:32]   = Image[822];
    assign  image_0_741[31:24]   = Image[823];
    assign  image_0_741[23:16]   = Image[853];
    assign  image_0_741[15:8]    = Image[854];
    assign  image_0_741[7:0]     = Image[855];

    assign  image_0_742[71:64]   = Image[790];
    assign  image_0_742[63:56]   = Image[791];
    assign  image_0_742[55:48]   = Image[792];
    assign  image_0_742[47:40]   = Image[822];
    assign  image_0_742[39:32]   = Image[823];
    assign  image_0_742[31:24]   = Image[824];
    assign  image_0_742[23:16]   = Image[854];
    assign  image_0_742[15:8]    = Image[855];
    assign  image_0_742[7:0]     = Image[856];

    assign  image_0_743[71:64]   = Image[791];
    assign  image_0_743[63:56]   = Image[792];
    assign  image_0_743[55:48]   = Image[793];
    assign  image_0_743[47:40]   = Image[823];
    assign  image_0_743[39:32]   = Image[824];
    assign  image_0_743[31:24]   = Image[825];
    assign  image_0_743[23:16]   = Image[855];
    assign  image_0_743[15:8]    = Image[856];
    assign  image_0_743[7:0]     = Image[857];

    assign  image_0_744[71:64]   = Image[792];
    assign  image_0_744[63:56]   = Image[793];
    assign  image_0_744[55:48]   = Image[794];
    assign  image_0_744[47:40]   = Image[824];
    assign  image_0_744[39:32]   = Image[825];
    assign  image_0_744[31:24]   = Image[826];
    assign  image_0_744[23:16]   = Image[856];
    assign  image_0_744[15:8]    = Image[857];
    assign  image_0_744[7:0]     = Image[858];

    assign  image_0_745[71:64]   = Image[793];
    assign  image_0_745[63:56]   = Image[794];
    assign  image_0_745[55:48]   = Image[795];
    assign  image_0_745[47:40]   = Image[825];
    assign  image_0_745[39:32]   = Image[826];
    assign  image_0_745[31:24]   = Image[827];
    assign  image_0_745[23:16]   = Image[857];
    assign  image_0_745[15:8]    = Image[858];
    assign  image_0_745[7:0]     = Image[859];

    assign  image_0_746[71:64]   = Image[794];
    assign  image_0_746[63:56]   = Image[795];
    assign  image_0_746[55:48]   = Image[796];
    assign  image_0_746[47:40]   = Image[826];
    assign  image_0_746[39:32]   = Image[827];
    assign  image_0_746[31:24]   = Image[828];
    assign  image_0_746[23:16]   = Image[858];
    assign  image_0_746[15:8]    = Image[859];
    assign  image_0_746[7:0]     = Image[860];

    assign  image_0_747[71:64]   = Image[795];
    assign  image_0_747[63:56]   = Image[796];
    assign  image_0_747[55:48]   = Image[797];
    assign  image_0_747[47:40]   = Image[827];
    assign  image_0_747[39:32]   = Image[828];
    assign  image_0_747[31:24]   = Image[829];
    assign  image_0_747[23:16]   = Image[859];
    assign  image_0_747[15:8]    = Image[860];
    assign  image_0_747[7:0]     = Image[861];

    assign  image_0_748[71:64]   = Image[796];
    assign  image_0_748[63:56]   = Image[797];
    assign  image_0_748[55:48]   = Image[798];
    assign  image_0_748[47:40]   = Image[828];
    assign  image_0_748[39:32]   = Image[829];
    assign  image_0_748[31:24]   = Image[830];
    assign  image_0_748[23:16]   = Image[860];
    assign  image_0_748[15:8]    = Image[861];
    assign  image_0_748[7:0]     = Image[862];

    assign  image_0_749[71:64]   = Image[797];
    assign  image_0_749[63:56]   = Image[798];
    assign  image_0_749[55:48]   = Image[799];
    assign  image_0_749[47:40]   = Image[829];
    assign  image_0_749[39:32]   = Image[830];
    assign  image_0_749[31:24]   = Image[831];
    assign  image_0_749[23:16]   = Image[861];
    assign  image_0_749[15:8]    = Image[862];
    assign  image_0_749[7:0]     = Image[863];

    assign  image_0_750[71:64]   = Image[800];
    assign  image_0_750[63:56]   = Image[801];
    assign  image_0_750[55:48]   = Image[802];
    assign  image_0_750[47:40]   = Image[832];
    assign  image_0_750[39:32]   = Image[833];
    assign  image_0_750[31:24]   = Image[834];
    assign  image_0_750[23:16]   = Image[864];
    assign  image_0_750[15:8]    = Image[865];
    assign  image_0_750[7:0]     = Image[866];

    assign  image_0_751[71:64]   = Image[801];
    assign  image_0_751[63:56]   = Image[802];
    assign  image_0_751[55:48]   = Image[803];
    assign  image_0_751[47:40]   = Image[833];
    assign  image_0_751[39:32]   = Image[834];
    assign  image_0_751[31:24]   = Image[835];
    assign  image_0_751[23:16]   = Image[865];
    assign  image_0_751[15:8]    = Image[866];
    assign  image_0_751[7:0]     = Image[867];

    assign  image_0_752[71:64]   = Image[802];
    assign  image_0_752[63:56]   = Image[803];
    assign  image_0_752[55:48]   = Image[804];
    assign  image_0_752[47:40]   = Image[834];
    assign  image_0_752[39:32]   = Image[835];
    assign  image_0_752[31:24]   = Image[836];
    assign  image_0_752[23:16]   = Image[866];
    assign  image_0_752[15:8]    = Image[867];
    assign  image_0_752[7:0]     = Image[868];

    assign  image_0_753[71:64]   = Image[803];
    assign  image_0_753[63:56]   = Image[804];
    assign  image_0_753[55:48]   = Image[805];
    assign  image_0_753[47:40]   = Image[835];
    assign  image_0_753[39:32]   = Image[836];
    assign  image_0_753[31:24]   = Image[837];
    assign  image_0_753[23:16]   = Image[867];
    assign  image_0_753[15:8]    = Image[868];
    assign  image_0_753[7:0]     = Image[869];

    assign  image_0_754[71:64]   = Image[804];
    assign  image_0_754[63:56]   = Image[805];
    assign  image_0_754[55:48]   = Image[806];
    assign  image_0_754[47:40]   = Image[836];
    assign  image_0_754[39:32]   = Image[837];
    assign  image_0_754[31:24]   = Image[838];
    assign  image_0_754[23:16]   = Image[868];
    assign  image_0_754[15:8]    = Image[869];
    assign  image_0_754[7:0]     = Image[870];

    assign  image_0_755[71:64]   = Image[805];
    assign  image_0_755[63:56]   = Image[806];
    assign  image_0_755[55:48]   = Image[807];
    assign  image_0_755[47:40]   = Image[837];
    assign  image_0_755[39:32]   = Image[838];
    assign  image_0_755[31:24]   = Image[839];
    assign  image_0_755[23:16]   = Image[869];
    assign  image_0_755[15:8]    = Image[870];
    assign  image_0_755[7:0]     = Image[871];

    assign  image_0_756[71:64]   = Image[806];
    assign  image_0_756[63:56]   = Image[807];
    assign  image_0_756[55:48]   = Image[808];
    assign  image_0_756[47:40]   = Image[838];
    assign  image_0_756[39:32]   = Image[839];
    assign  image_0_756[31:24]   = Image[840];
    assign  image_0_756[23:16]   = Image[870];
    assign  image_0_756[15:8]    = Image[871];
    assign  image_0_756[7:0]     = Image[872];

    assign  image_0_757[71:64]   = Image[807];
    assign  image_0_757[63:56]   = Image[808];
    assign  image_0_757[55:48]   = Image[809];
    assign  image_0_757[47:40]   = Image[839];
    assign  image_0_757[39:32]   = Image[840];
    assign  image_0_757[31:24]   = Image[841];
    assign  image_0_757[23:16]   = Image[871];
    assign  image_0_757[15:8]    = Image[872];
    assign  image_0_757[7:0]     = Image[873];

    assign  image_0_758[71:64]   = Image[808];
    assign  image_0_758[63:56]   = Image[809];
    assign  image_0_758[55:48]   = Image[810];
    assign  image_0_758[47:40]   = Image[840];
    assign  image_0_758[39:32]   = Image[841];
    assign  image_0_758[31:24]   = Image[842];
    assign  image_0_758[23:16]   = Image[872];
    assign  image_0_758[15:8]    = Image[873];
    assign  image_0_758[7:0]     = Image[874];

    assign  image_0_759[71:64]   = Image[809];
    assign  image_0_759[63:56]   = Image[810];
    assign  image_0_759[55:48]   = Image[811];
    assign  image_0_759[47:40]   = Image[841];
    assign  image_0_759[39:32]   = Image[842];
    assign  image_0_759[31:24]   = Image[843];
    assign  image_0_759[23:16]   = Image[873];
    assign  image_0_759[15:8]    = Image[874];
    assign  image_0_759[7:0]     = Image[875];

    assign  image_0_760[71:64]   = Image[810];
    assign  image_0_760[63:56]   = Image[811];
    assign  image_0_760[55:48]   = Image[812];
    assign  image_0_760[47:40]   = Image[842];
    assign  image_0_760[39:32]   = Image[843];
    assign  image_0_760[31:24]   = Image[844];
    assign  image_0_760[23:16]   = Image[874];
    assign  image_0_760[15:8]    = Image[875];
    assign  image_0_760[7:0]     = Image[876];

    assign  image_0_761[71:64]   = Image[811];
    assign  image_0_761[63:56]   = Image[812];
    assign  image_0_761[55:48]   = Image[813];
    assign  image_0_761[47:40]   = Image[843];
    assign  image_0_761[39:32]   = Image[844];
    assign  image_0_761[31:24]   = Image[845];
    assign  image_0_761[23:16]   = Image[875];
    assign  image_0_761[15:8]    = Image[876];
    assign  image_0_761[7:0]     = Image[877];

    assign  image_0_762[71:64]   = Image[812];
    assign  image_0_762[63:56]   = Image[813];
    assign  image_0_762[55:48]   = Image[814];
    assign  image_0_762[47:40]   = Image[844];
    assign  image_0_762[39:32]   = Image[845];
    assign  image_0_762[31:24]   = Image[846];
    assign  image_0_762[23:16]   = Image[876];
    assign  image_0_762[15:8]    = Image[877];
    assign  image_0_762[7:0]     = Image[878];

    assign  image_0_763[71:64]   = Image[813];
    assign  image_0_763[63:56]   = Image[814];
    assign  image_0_763[55:48]   = Image[815];
    assign  image_0_763[47:40]   = Image[845];
    assign  image_0_763[39:32]   = Image[846];
    assign  image_0_763[31:24]   = Image[847];
    assign  image_0_763[23:16]   = Image[877];
    assign  image_0_763[15:8]    = Image[878];
    assign  image_0_763[7:0]     = Image[879];

    assign  image_0_764[71:64]   = Image[814];
    assign  image_0_764[63:56]   = Image[815];
    assign  image_0_764[55:48]   = Image[816];
    assign  image_0_764[47:40]   = Image[846];
    assign  image_0_764[39:32]   = Image[847];
    assign  image_0_764[31:24]   = Image[848];
    assign  image_0_764[23:16]   = Image[878];
    assign  image_0_764[15:8]    = Image[879];
    assign  image_0_764[7:0]     = Image[880];

    assign  image_0_765[71:64]   = Image[815];
    assign  image_0_765[63:56]   = Image[816];
    assign  image_0_765[55:48]   = Image[817];
    assign  image_0_765[47:40]   = Image[847];
    assign  image_0_765[39:32]   = Image[848];
    assign  image_0_765[31:24]   = Image[849];
    assign  image_0_765[23:16]   = Image[879];
    assign  image_0_765[15:8]    = Image[880];
    assign  image_0_765[7:0]     = Image[881];

    assign  image_0_766[71:64]   = Image[816];
    assign  image_0_766[63:56]   = Image[817];
    assign  image_0_766[55:48]   = Image[818];
    assign  image_0_766[47:40]   = Image[848];
    assign  image_0_766[39:32]   = Image[849];
    assign  image_0_766[31:24]   = Image[850];
    assign  image_0_766[23:16]   = Image[880];
    assign  image_0_766[15:8]    = Image[881];
    assign  image_0_766[7:0]     = Image[882];

    assign  image_0_767[71:64]   = Image[817];
    assign  image_0_767[63:56]   = Image[818];
    assign  image_0_767[55:48]   = Image[819];
    assign  image_0_767[47:40]   = Image[849];
    assign  image_0_767[39:32]   = Image[850];
    assign  image_0_767[31:24]   = Image[851];
    assign  image_0_767[23:16]   = Image[881];
    assign  image_0_767[15:8]    = Image[882];
    assign  image_0_767[7:0]     = Image[883];

    assign  image_0_768[71:64]   = Image[818];
    assign  image_0_768[63:56]   = Image[819];
    assign  image_0_768[55:48]   = Image[820];
    assign  image_0_768[47:40]   = Image[850];
    assign  image_0_768[39:32]   = Image[851];
    assign  image_0_768[31:24]   = Image[852];
    assign  image_0_768[23:16]   = Image[882];
    assign  image_0_768[15:8]    = Image[883];
    assign  image_0_768[7:0]     = Image[884];

    assign  image_0_769[71:64]   = Image[819];
    assign  image_0_769[63:56]   = Image[820];
    assign  image_0_769[55:48]   = Image[821];
    assign  image_0_769[47:40]   = Image[851];
    assign  image_0_769[39:32]   = Image[852];
    assign  image_0_769[31:24]   = Image[853];
    assign  image_0_769[23:16]   = Image[883];
    assign  image_0_769[15:8]    = Image[884];
    assign  image_0_769[7:0]     = Image[885];

    assign  image_0_770[71:64]   = Image[820];
    assign  image_0_770[63:56]   = Image[821];
    assign  image_0_770[55:48]   = Image[822];
    assign  image_0_770[47:40]   = Image[852];
    assign  image_0_770[39:32]   = Image[853];
    assign  image_0_770[31:24]   = Image[854];
    assign  image_0_770[23:16]   = Image[884];
    assign  image_0_770[15:8]    = Image[885];
    assign  image_0_770[7:0]     = Image[886];

    assign  image_0_771[71:64]   = Image[821];
    assign  image_0_771[63:56]   = Image[822];
    assign  image_0_771[55:48]   = Image[823];
    assign  image_0_771[47:40]   = Image[853];
    assign  image_0_771[39:32]   = Image[854];
    assign  image_0_771[31:24]   = Image[855];
    assign  image_0_771[23:16]   = Image[885];
    assign  image_0_771[15:8]    = Image[886];
    assign  image_0_771[7:0]     = Image[887];

    assign  image_0_772[71:64]   = Image[822];
    assign  image_0_772[63:56]   = Image[823];
    assign  image_0_772[55:48]   = Image[824];
    assign  image_0_772[47:40]   = Image[854];
    assign  image_0_772[39:32]   = Image[855];
    assign  image_0_772[31:24]   = Image[856];
    assign  image_0_772[23:16]   = Image[886];
    assign  image_0_772[15:8]    = Image[887];
    assign  image_0_772[7:0]     = Image[888];

    assign  image_0_773[71:64]   = Image[823];
    assign  image_0_773[63:56]   = Image[824];
    assign  image_0_773[55:48]   = Image[825];
    assign  image_0_773[47:40]   = Image[855];
    assign  image_0_773[39:32]   = Image[856];
    assign  image_0_773[31:24]   = Image[857];
    assign  image_0_773[23:16]   = Image[887];
    assign  image_0_773[15:8]    = Image[888];
    assign  image_0_773[7:0]     = Image[889];

    assign  image_0_774[71:64]   = Image[824];
    assign  image_0_774[63:56]   = Image[825];
    assign  image_0_774[55:48]   = Image[826];
    assign  image_0_774[47:40]   = Image[856];
    assign  image_0_774[39:32]   = Image[857];
    assign  image_0_774[31:24]   = Image[858];
    assign  image_0_774[23:16]   = Image[888];
    assign  image_0_774[15:8]    = Image[889];
    assign  image_0_774[7:0]     = Image[890];

    assign  image_0_775[71:64]   = Image[825];
    assign  image_0_775[63:56]   = Image[826];
    assign  image_0_775[55:48]   = Image[827];
    assign  image_0_775[47:40]   = Image[857];
    assign  image_0_775[39:32]   = Image[858];
    assign  image_0_775[31:24]   = Image[859];
    assign  image_0_775[23:16]   = Image[889];
    assign  image_0_775[15:8]    = Image[890];
    assign  image_0_775[7:0]     = Image[891];

    assign  image_0_776[71:64]   = Image[826];
    assign  image_0_776[63:56]   = Image[827];
    assign  image_0_776[55:48]   = Image[828];
    assign  image_0_776[47:40]   = Image[858];
    assign  image_0_776[39:32]   = Image[859];
    assign  image_0_776[31:24]   = Image[860];
    assign  image_0_776[23:16]   = Image[890];
    assign  image_0_776[15:8]    = Image[891];
    assign  image_0_776[7:0]     = Image[892];

    assign  image_0_777[71:64]   = Image[827];
    assign  image_0_777[63:56]   = Image[828];
    assign  image_0_777[55:48]   = Image[829];
    assign  image_0_777[47:40]   = Image[859];
    assign  image_0_777[39:32]   = Image[860];
    assign  image_0_777[31:24]   = Image[861];
    assign  image_0_777[23:16]   = Image[891];
    assign  image_0_777[15:8]    = Image[892];
    assign  image_0_777[7:0]     = Image[893];

    assign  image_0_778[71:64]   = Image[828];
    assign  image_0_778[63:56]   = Image[829];
    assign  image_0_778[55:48]   = Image[830];
    assign  image_0_778[47:40]   = Image[860];
    assign  image_0_778[39:32]   = Image[861];
    assign  image_0_778[31:24]   = Image[862];
    assign  image_0_778[23:16]   = Image[892];
    assign  image_0_778[15:8]    = Image[893];
    assign  image_0_778[7:0]     = Image[894];

    assign  image_0_779[71:64]   = Image[829];
    assign  image_0_779[63:56]   = Image[830];
    assign  image_0_779[55:48]   = Image[831];
    assign  image_0_779[47:40]   = Image[861];
    assign  image_0_779[39:32]   = Image[862];
    assign  image_0_779[31:24]   = Image[863];
    assign  image_0_779[23:16]   = Image[893];
    assign  image_0_779[15:8]    = Image[894];
    assign  image_0_779[7:0]     = Image[895];

    assign  image_0_780[71:64]   = Image[832];
    assign  image_0_780[63:56]   = Image[833];
    assign  image_0_780[55:48]   = Image[834];
    assign  image_0_780[47:40]   = Image[864];
    assign  image_0_780[39:32]   = Image[865];
    assign  image_0_780[31:24]   = Image[866];
    assign  image_0_780[23:16]   = Image[896];
    assign  image_0_780[15:8]    = Image[897];
    assign  image_0_780[7:0]     = Image[898];

    assign  image_0_781[71:64]   = Image[833];
    assign  image_0_781[63:56]   = Image[834];
    assign  image_0_781[55:48]   = Image[835];
    assign  image_0_781[47:40]   = Image[865];
    assign  image_0_781[39:32]   = Image[866];
    assign  image_0_781[31:24]   = Image[867];
    assign  image_0_781[23:16]   = Image[897];
    assign  image_0_781[15:8]    = Image[898];
    assign  image_0_781[7:0]     = Image[899];

    assign  image_0_782[71:64]   = Image[834];
    assign  image_0_782[63:56]   = Image[835];
    assign  image_0_782[55:48]   = Image[836];
    assign  image_0_782[47:40]   = Image[866];
    assign  image_0_782[39:32]   = Image[867];
    assign  image_0_782[31:24]   = Image[868];
    assign  image_0_782[23:16]   = Image[898];
    assign  image_0_782[15:8]    = Image[899];
    assign  image_0_782[7:0]     = Image[900];

    assign  image_0_783[71:64]   = Image[835];
    assign  image_0_783[63:56]   = Image[836];
    assign  image_0_783[55:48]   = Image[837];
    assign  image_0_783[47:40]   = Image[867];
    assign  image_0_783[39:32]   = Image[868];
    assign  image_0_783[31:24]   = Image[869];
    assign  image_0_783[23:16]   = Image[899];
    assign  image_0_783[15:8]    = Image[900];
    assign  image_0_783[7:0]     = Image[901];

    assign  image_0_784[71:64]   = Image[836];
    assign  image_0_784[63:56]   = Image[837];
    assign  image_0_784[55:48]   = Image[838];
    assign  image_0_784[47:40]   = Image[868];
    assign  image_0_784[39:32]   = Image[869];
    assign  image_0_784[31:24]   = Image[870];
    assign  image_0_784[23:16]   = Image[900];
    assign  image_0_784[15:8]    = Image[901];
    assign  image_0_784[7:0]     = Image[902];

    assign  image_0_785[71:64]   = Image[837];
    assign  image_0_785[63:56]   = Image[838];
    assign  image_0_785[55:48]   = Image[839];
    assign  image_0_785[47:40]   = Image[869];
    assign  image_0_785[39:32]   = Image[870];
    assign  image_0_785[31:24]   = Image[871];
    assign  image_0_785[23:16]   = Image[901];
    assign  image_0_785[15:8]    = Image[902];
    assign  image_0_785[7:0]     = Image[903];

    assign  image_0_786[71:64]   = Image[838];
    assign  image_0_786[63:56]   = Image[839];
    assign  image_0_786[55:48]   = Image[840];
    assign  image_0_786[47:40]   = Image[870];
    assign  image_0_786[39:32]   = Image[871];
    assign  image_0_786[31:24]   = Image[872];
    assign  image_0_786[23:16]   = Image[902];
    assign  image_0_786[15:8]    = Image[903];
    assign  image_0_786[7:0]     = Image[904];

    assign  image_0_787[71:64]   = Image[839];
    assign  image_0_787[63:56]   = Image[840];
    assign  image_0_787[55:48]   = Image[841];
    assign  image_0_787[47:40]   = Image[871];
    assign  image_0_787[39:32]   = Image[872];
    assign  image_0_787[31:24]   = Image[873];
    assign  image_0_787[23:16]   = Image[903];
    assign  image_0_787[15:8]    = Image[904];
    assign  image_0_787[7:0]     = Image[905];

    assign  image_0_788[71:64]   = Image[840];
    assign  image_0_788[63:56]   = Image[841];
    assign  image_0_788[55:48]   = Image[842];
    assign  image_0_788[47:40]   = Image[872];
    assign  image_0_788[39:32]   = Image[873];
    assign  image_0_788[31:24]   = Image[874];
    assign  image_0_788[23:16]   = Image[904];
    assign  image_0_788[15:8]    = Image[905];
    assign  image_0_788[7:0]     = Image[906];

    assign  image_0_789[71:64]   = Image[841];
    assign  image_0_789[63:56]   = Image[842];
    assign  image_0_789[55:48]   = Image[843];
    assign  image_0_789[47:40]   = Image[873];
    assign  image_0_789[39:32]   = Image[874];
    assign  image_0_789[31:24]   = Image[875];
    assign  image_0_789[23:16]   = Image[905];
    assign  image_0_789[15:8]    = Image[906];
    assign  image_0_789[7:0]     = Image[907];

    assign  image_0_790[71:64]   = Image[842];
    assign  image_0_790[63:56]   = Image[843];
    assign  image_0_790[55:48]   = Image[844];
    assign  image_0_790[47:40]   = Image[874];
    assign  image_0_790[39:32]   = Image[875];
    assign  image_0_790[31:24]   = Image[876];
    assign  image_0_790[23:16]   = Image[906];
    assign  image_0_790[15:8]    = Image[907];
    assign  image_0_790[7:0]     = Image[908];

    assign  image_0_791[71:64]   = Image[843];
    assign  image_0_791[63:56]   = Image[844];
    assign  image_0_791[55:48]   = Image[845];
    assign  image_0_791[47:40]   = Image[875];
    assign  image_0_791[39:32]   = Image[876];
    assign  image_0_791[31:24]   = Image[877];
    assign  image_0_791[23:16]   = Image[907];
    assign  image_0_791[15:8]    = Image[908];
    assign  image_0_791[7:0]     = Image[909];

    assign  image_0_792[71:64]   = Image[844];
    assign  image_0_792[63:56]   = Image[845];
    assign  image_0_792[55:48]   = Image[846];
    assign  image_0_792[47:40]   = Image[876];
    assign  image_0_792[39:32]   = Image[877];
    assign  image_0_792[31:24]   = Image[878];
    assign  image_0_792[23:16]   = Image[908];
    assign  image_0_792[15:8]    = Image[909];
    assign  image_0_792[7:0]     = Image[910];

    assign  image_0_793[71:64]   = Image[845];
    assign  image_0_793[63:56]   = Image[846];
    assign  image_0_793[55:48]   = Image[847];
    assign  image_0_793[47:40]   = Image[877];
    assign  image_0_793[39:32]   = Image[878];
    assign  image_0_793[31:24]   = Image[879];
    assign  image_0_793[23:16]   = Image[909];
    assign  image_0_793[15:8]    = Image[910];
    assign  image_0_793[7:0]     = Image[911];

    assign  image_0_794[71:64]   = Image[846];
    assign  image_0_794[63:56]   = Image[847];
    assign  image_0_794[55:48]   = Image[848];
    assign  image_0_794[47:40]   = Image[878];
    assign  image_0_794[39:32]   = Image[879];
    assign  image_0_794[31:24]   = Image[880];
    assign  image_0_794[23:16]   = Image[910];
    assign  image_0_794[15:8]    = Image[911];
    assign  image_0_794[7:0]     = Image[912];

    assign  image_0_795[71:64]   = Image[847];
    assign  image_0_795[63:56]   = Image[848];
    assign  image_0_795[55:48]   = Image[849];
    assign  image_0_795[47:40]   = Image[879];
    assign  image_0_795[39:32]   = Image[880];
    assign  image_0_795[31:24]   = Image[881];
    assign  image_0_795[23:16]   = Image[911];
    assign  image_0_795[15:8]    = Image[912];
    assign  image_0_795[7:0]     = Image[913];

    assign  image_0_796[71:64]   = Image[848];
    assign  image_0_796[63:56]   = Image[849];
    assign  image_0_796[55:48]   = Image[850];
    assign  image_0_796[47:40]   = Image[880];
    assign  image_0_796[39:32]   = Image[881];
    assign  image_0_796[31:24]   = Image[882];
    assign  image_0_796[23:16]   = Image[912];
    assign  image_0_796[15:8]    = Image[913];
    assign  image_0_796[7:0]     = Image[914];

    assign  image_0_797[71:64]   = Image[849];
    assign  image_0_797[63:56]   = Image[850];
    assign  image_0_797[55:48]   = Image[851];
    assign  image_0_797[47:40]   = Image[881];
    assign  image_0_797[39:32]   = Image[882];
    assign  image_0_797[31:24]   = Image[883];
    assign  image_0_797[23:16]   = Image[913];
    assign  image_0_797[15:8]    = Image[914];
    assign  image_0_797[7:0]     = Image[915];

    assign  image_0_798[71:64]   = Image[850];
    assign  image_0_798[63:56]   = Image[851];
    assign  image_0_798[55:48]   = Image[852];
    assign  image_0_798[47:40]   = Image[882];
    assign  image_0_798[39:32]   = Image[883];
    assign  image_0_798[31:24]   = Image[884];
    assign  image_0_798[23:16]   = Image[914];
    assign  image_0_798[15:8]    = Image[915];
    assign  image_0_798[7:0]     = Image[916];

    assign  image_0_799[71:64]   = Image[851];
    assign  image_0_799[63:56]   = Image[852];
    assign  image_0_799[55:48]   = Image[853];
    assign  image_0_799[47:40]   = Image[883];
    assign  image_0_799[39:32]   = Image[884];
    assign  image_0_799[31:24]   = Image[885];
    assign  image_0_799[23:16]   = Image[915];
    assign  image_0_799[15:8]    = Image[916];
    assign  image_0_799[7:0]     = Image[917];

    assign  image_0_800[71:64]   = Image[852];
    assign  image_0_800[63:56]   = Image[853];
    assign  image_0_800[55:48]   = Image[854];
    assign  image_0_800[47:40]   = Image[884];
    assign  image_0_800[39:32]   = Image[885];
    assign  image_0_800[31:24]   = Image[886];
    assign  image_0_800[23:16]   = Image[916];
    assign  image_0_800[15:8]    = Image[917];
    assign  image_0_800[7:0]     = Image[918];

    assign  image_0_801[71:64]   = Image[853];
    assign  image_0_801[63:56]   = Image[854];
    assign  image_0_801[55:48]   = Image[855];
    assign  image_0_801[47:40]   = Image[885];
    assign  image_0_801[39:32]   = Image[886];
    assign  image_0_801[31:24]   = Image[887];
    assign  image_0_801[23:16]   = Image[917];
    assign  image_0_801[15:8]    = Image[918];
    assign  image_0_801[7:0]     = Image[919];

    assign  image_0_802[71:64]   = Image[854];
    assign  image_0_802[63:56]   = Image[855];
    assign  image_0_802[55:48]   = Image[856];
    assign  image_0_802[47:40]   = Image[886];
    assign  image_0_802[39:32]   = Image[887];
    assign  image_0_802[31:24]   = Image[888];
    assign  image_0_802[23:16]   = Image[918];
    assign  image_0_802[15:8]    = Image[919];
    assign  image_0_802[7:0]     = Image[920];

    assign  image_0_803[71:64]   = Image[855];
    assign  image_0_803[63:56]   = Image[856];
    assign  image_0_803[55:48]   = Image[857];
    assign  image_0_803[47:40]   = Image[887];
    assign  image_0_803[39:32]   = Image[888];
    assign  image_0_803[31:24]   = Image[889];
    assign  image_0_803[23:16]   = Image[919];
    assign  image_0_803[15:8]    = Image[920];
    assign  image_0_803[7:0]     = Image[921];

    assign  image_0_804[71:64]   = Image[856];
    assign  image_0_804[63:56]   = Image[857];
    assign  image_0_804[55:48]   = Image[858];
    assign  image_0_804[47:40]   = Image[888];
    assign  image_0_804[39:32]   = Image[889];
    assign  image_0_804[31:24]   = Image[890];
    assign  image_0_804[23:16]   = Image[920];
    assign  image_0_804[15:8]    = Image[921];
    assign  image_0_804[7:0]     = Image[922];

    assign  image_0_805[71:64]   = Image[857];
    assign  image_0_805[63:56]   = Image[858];
    assign  image_0_805[55:48]   = Image[859];
    assign  image_0_805[47:40]   = Image[889];
    assign  image_0_805[39:32]   = Image[890];
    assign  image_0_805[31:24]   = Image[891];
    assign  image_0_805[23:16]   = Image[921];
    assign  image_0_805[15:8]    = Image[922];
    assign  image_0_805[7:0]     = Image[923];

    assign  image_0_806[71:64]   = Image[858];
    assign  image_0_806[63:56]   = Image[859];
    assign  image_0_806[55:48]   = Image[860];
    assign  image_0_806[47:40]   = Image[890];
    assign  image_0_806[39:32]   = Image[891];
    assign  image_0_806[31:24]   = Image[892];
    assign  image_0_806[23:16]   = Image[922];
    assign  image_0_806[15:8]    = Image[923];
    assign  image_0_806[7:0]     = Image[924];

    assign  image_0_807[71:64]   = Image[859];
    assign  image_0_807[63:56]   = Image[860];
    assign  image_0_807[55:48]   = Image[861];
    assign  image_0_807[47:40]   = Image[891];
    assign  image_0_807[39:32]   = Image[892];
    assign  image_0_807[31:24]   = Image[893];
    assign  image_0_807[23:16]   = Image[923];
    assign  image_0_807[15:8]    = Image[924];
    assign  image_0_807[7:0]     = Image[925];

    assign  image_0_808[71:64]   = Image[860];
    assign  image_0_808[63:56]   = Image[861];
    assign  image_0_808[55:48]   = Image[862];
    assign  image_0_808[47:40]   = Image[892];
    assign  image_0_808[39:32]   = Image[893];
    assign  image_0_808[31:24]   = Image[894];
    assign  image_0_808[23:16]   = Image[924];
    assign  image_0_808[15:8]    = Image[925];
    assign  image_0_808[7:0]     = Image[926];

    assign  image_0_809[71:64]   = Image[861];
    assign  image_0_809[63:56]   = Image[862];
    assign  image_0_809[55:48]   = Image[863];
    assign  image_0_809[47:40]   = Image[893];
    assign  image_0_809[39:32]   = Image[894];
    assign  image_0_809[31:24]   = Image[895];
    assign  image_0_809[23:16]   = Image[925];
    assign  image_0_809[15:8]    = Image[926];
    assign  image_0_809[7:0]     = Image[927];

    assign  image_0_810[71:64]   = Image[864];
    assign  image_0_810[63:56]   = Image[865];
    assign  image_0_810[55:48]   = Image[866];
    assign  image_0_810[47:40]   = Image[896];
    assign  image_0_810[39:32]   = Image[897];
    assign  image_0_810[31:24]   = Image[898];
    assign  image_0_810[23:16]   = Image[928];
    assign  image_0_810[15:8]    = Image[929];
    assign  image_0_810[7:0]     = Image[930];

    assign  image_0_811[71:64]   = Image[865];
    assign  image_0_811[63:56]   = Image[866];
    assign  image_0_811[55:48]   = Image[867];
    assign  image_0_811[47:40]   = Image[897];
    assign  image_0_811[39:32]   = Image[898];
    assign  image_0_811[31:24]   = Image[899];
    assign  image_0_811[23:16]   = Image[929];
    assign  image_0_811[15:8]    = Image[930];
    assign  image_0_811[7:0]     = Image[931];

    assign  image_0_812[71:64]   = Image[866];
    assign  image_0_812[63:56]   = Image[867];
    assign  image_0_812[55:48]   = Image[868];
    assign  image_0_812[47:40]   = Image[898];
    assign  image_0_812[39:32]   = Image[899];
    assign  image_0_812[31:24]   = Image[900];
    assign  image_0_812[23:16]   = Image[930];
    assign  image_0_812[15:8]    = Image[931];
    assign  image_0_812[7:0]     = Image[932];

    assign  image_0_813[71:64]   = Image[867];
    assign  image_0_813[63:56]   = Image[868];
    assign  image_0_813[55:48]   = Image[869];
    assign  image_0_813[47:40]   = Image[899];
    assign  image_0_813[39:32]   = Image[900];
    assign  image_0_813[31:24]   = Image[901];
    assign  image_0_813[23:16]   = Image[931];
    assign  image_0_813[15:8]    = Image[932];
    assign  image_0_813[7:0]     = Image[933];

    assign  image_0_814[71:64]   = Image[868];
    assign  image_0_814[63:56]   = Image[869];
    assign  image_0_814[55:48]   = Image[870];
    assign  image_0_814[47:40]   = Image[900];
    assign  image_0_814[39:32]   = Image[901];
    assign  image_0_814[31:24]   = Image[902];
    assign  image_0_814[23:16]   = Image[932];
    assign  image_0_814[15:8]    = Image[933];
    assign  image_0_814[7:0]     = Image[934];

    assign  image_0_815[71:64]   = Image[869];
    assign  image_0_815[63:56]   = Image[870];
    assign  image_0_815[55:48]   = Image[871];
    assign  image_0_815[47:40]   = Image[901];
    assign  image_0_815[39:32]   = Image[902];
    assign  image_0_815[31:24]   = Image[903];
    assign  image_0_815[23:16]   = Image[933];
    assign  image_0_815[15:8]    = Image[934];
    assign  image_0_815[7:0]     = Image[935];

    assign  image_0_816[71:64]   = Image[870];
    assign  image_0_816[63:56]   = Image[871];
    assign  image_0_816[55:48]   = Image[872];
    assign  image_0_816[47:40]   = Image[902];
    assign  image_0_816[39:32]   = Image[903];
    assign  image_0_816[31:24]   = Image[904];
    assign  image_0_816[23:16]   = Image[934];
    assign  image_0_816[15:8]    = Image[935];
    assign  image_0_816[7:0]     = Image[936];

    assign  image_0_817[71:64]   = Image[871];
    assign  image_0_817[63:56]   = Image[872];
    assign  image_0_817[55:48]   = Image[873];
    assign  image_0_817[47:40]   = Image[903];
    assign  image_0_817[39:32]   = Image[904];
    assign  image_0_817[31:24]   = Image[905];
    assign  image_0_817[23:16]   = Image[935];
    assign  image_0_817[15:8]    = Image[936];
    assign  image_0_817[7:0]     = Image[937];

    assign  image_0_818[71:64]   = Image[872];
    assign  image_0_818[63:56]   = Image[873];
    assign  image_0_818[55:48]   = Image[874];
    assign  image_0_818[47:40]   = Image[904];
    assign  image_0_818[39:32]   = Image[905];
    assign  image_0_818[31:24]   = Image[906];
    assign  image_0_818[23:16]   = Image[936];
    assign  image_0_818[15:8]    = Image[937];
    assign  image_0_818[7:0]     = Image[938];

    assign  image_0_819[71:64]   = Image[873];
    assign  image_0_819[63:56]   = Image[874];
    assign  image_0_819[55:48]   = Image[875];
    assign  image_0_819[47:40]   = Image[905];
    assign  image_0_819[39:32]   = Image[906];
    assign  image_0_819[31:24]   = Image[907];
    assign  image_0_819[23:16]   = Image[937];
    assign  image_0_819[15:8]    = Image[938];
    assign  image_0_819[7:0]     = Image[939];

    assign  image_0_820[71:64]   = Image[874];
    assign  image_0_820[63:56]   = Image[875];
    assign  image_0_820[55:48]   = Image[876];
    assign  image_0_820[47:40]   = Image[906];
    assign  image_0_820[39:32]   = Image[907];
    assign  image_0_820[31:24]   = Image[908];
    assign  image_0_820[23:16]   = Image[938];
    assign  image_0_820[15:8]    = Image[939];
    assign  image_0_820[7:0]     = Image[940];

    assign  image_0_821[71:64]   = Image[875];
    assign  image_0_821[63:56]   = Image[876];
    assign  image_0_821[55:48]   = Image[877];
    assign  image_0_821[47:40]   = Image[907];
    assign  image_0_821[39:32]   = Image[908];
    assign  image_0_821[31:24]   = Image[909];
    assign  image_0_821[23:16]   = Image[939];
    assign  image_0_821[15:8]    = Image[940];
    assign  image_0_821[7:0]     = Image[941];

    assign  image_0_822[71:64]   = Image[876];
    assign  image_0_822[63:56]   = Image[877];
    assign  image_0_822[55:48]   = Image[878];
    assign  image_0_822[47:40]   = Image[908];
    assign  image_0_822[39:32]   = Image[909];
    assign  image_0_822[31:24]   = Image[910];
    assign  image_0_822[23:16]   = Image[940];
    assign  image_0_822[15:8]    = Image[941];
    assign  image_0_822[7:0]     = Image[942];

    assign  image_0_823[71:64]   = Image[877];
    assign  image_0_823[63:56]   = Image[878];
    assign  image_0_823[55:48]   = Image[879];
    assign  image_0_823[47:40]   = Image[909];
    assign  image_0_823[39:32]   = Image[910];
    assign  image_0_823[31:24]   = Image[911];
    assign  image_0_823[23:16]   = Image[941];
    assign  image_0_823[15:8]    = Image[942];
    assign  image_0_823[7:0]     = Image[943];

    assign  image_0_824[71:64]   = Image[878];
    assign  image_0_824[63:56]   = Image[879];
    assign  image_0_824[55:48]   = Image[880];
    assign  image_0_824[47:40]   = Image[910];
    assign  image_0_824[39:32]   = Image[911];
    assign  image_0_824[31:24]   = Image[912];
    assign  image_0_824[23:16]   = Image[942];
    assign  image_0_824[15:8]    = Image[943];
    assign  image_0_824[7:0]     = Image[944];

    assign  image_0_825[71:64]   = Image[879];
    assign  image_0_825[63:56]   = Image[880];
    assign  image_0_825[55:48]   = Image[881];
    assign  image_0_825[47:40]   = Image[911];
    assign  image_0_825[39:32]   = Image[912];
    assign  image_0_825[31:24]   = Image[913];
    assign  image_0_825[23:16]   = Image[943];
    assign  image_0_825[15:8]    = Image[944];
    assign  image_0_825[7:0]     = Image[945];

    assign  image_0_826[71:64]   = Image[880];
    assign  image_0_826[63:56]   = Image[881];
    assign  image_0_826[55:48]   = Image[882];
    assign  image_0_826[47:40]   = Image[912];
    assign  image_0_826[39:32]   = Image[913];
    assign  image_0_826[31:24]   = Image[914];
    assign  image_0_826[23:16]   = Image[944];
    assign  image_0_826[15:8]    = Image[945];
    assign  image_0_826[7:0]     = Image[946];

    assign  image_0_827[71:64]   = Image[881];
    assign  image_0_827[63:56]   = Image[882];
    assign  image_0_827[55:48]   = Image[883];
    assign  image_0_827[47:40]   = Image[913];
    assign  image_0_827[39:32]   = Image[914];
    assign  image_0_827[31:24]   = Image[915];
    assign  image_0_827[23:16]   = Image[945];
    assign  image_0_827[15:8]    = Image[946];
    assign  image_0_827[7:0]     = Image[947];

    assign  image_0_828[71:64]   = Image[882];
    assign  image_0_828[63:56]   = Image[883];
    assign  image_0_828[55:48]   = Image[884];
    assign  image_0_828[47:40]   = Image[914];
    assign  image_0_828[39:32]   = Image[915];
    assign  image_0_828[31:24]   = Image[916];
    assign  image_0_828[23:16]   = Image[946];
    assign  image_0_828[15:8]    = Image[947];
    assign  image_0_828[7:0]     = Image[948];

    assign  image_0_829[71:64]   = Image[883];
    assign  image_0_829[63:56]   = Image[884];
    assign  image_0_829[55:48]   = Image[885];
    assign  image_0_829[47:40]   = Image[915];
    assign  image_0_829[39:32]   = Image[916];
    assign  image_0_829[31:24]   = Image[917];
    assign  image_0_829[23:16]   = Image[947];
    assign  image_0_829[15:8]    = Image[948];
    assign  image_0_829[7:0]     = Image[949];

    assign  image_0_830[71:64]   = Image[884];
    assign  image_0_830[63:56]   = Image[885];
    assign  image_0_830[55:48]   = Image[886];
    assign  image_0_830[47:40]   = Image[916];
    assign  image_0_830[39:32]   = Image[917];
    assign  image_0_830[31:24]   = Image[918];
    assign  image_0_830[23:16]   = Image[948];
    assign  image_0_830[15:8]    = Image[949];
    assign  image_0_830[7:0]     = Image[950];

    assign  image_0_831[71:64]   = Image[885];
    assign  image_0_831[63:56]   = Image[886];
    assign  image_0_831[55:48]   = Image[887];
    assign  image_0_831[47:40]   = Image[917];
    assign  image_0_831[39:32]   = Image[918];
    assign  image_0_831[31:24]   = Image[919];
    assign  image_0_831[23:16]   = Image[949];
    assign  image_0_831[15:8]    = Image[950];
    assign  image_0_831[7:0]     = Image[951];

    assign  image_0_832[71:64]   = Image[886];
    assign  image_0_832[63:56]   = Image[887];
    assign  image_0_832[55:48]   = Image[888];
    assign  image_0_832[47:40]   = Image[918];
    assign  image_0_832[39:32]   = Image[919];
    assign  image_0_832[31:24]   = Image[920];
    assign  image_0_832[23:16]   = Image[950];
    assign  image_0_832[15:8]    = Image[951];
    assign  image_0_832[7:0]     = Image[952];

    assign  image_0_833[71:64]   = Image[887];
    assign  image_0_833[63:56]   = Image[888];
    assign  image_0_833[55:48]   = Image[889];
    assign  image_0_833[47:40]   = Image[919];
    assign  image_0_833[39:32]   = Image[920];
    assign  image_0_833[31:24]   = Image[921];
    assign  image_0_833[23:16]   = Image[951];
    assign  image_0_833[15:8]    = Image[952];
    assign  image_0_833[7:0]     = Image[953];

    assign  image_0_834[71:64]   = Image[888];
    assign  image_0_834[63:56]   = Image[889];
    assign  image_0_834[55:48]   = Image[890];
    assign  image_0_834[47:40]   = Image[920];
    assign  image_0_834[39:32]   = Image[921];
    assign  image_0_834[31:24]   = Image[922];
    assign  image_0_834[23:16]   = Image[952];
    assign  image_0_834[15:8]    = Image[953];
    assign  image_0_834[7:0]     = Image[954];

    assign  image_0_835[71:64]   = Image[889];
    assign  image_0_835[63:56]   = Image[890];
    assign  image_0_835[55:48]   = Image[891];
    assign  image_0_835[47:40]   = Image[921];
    assign  image_0_835[39:32]   = Image[922];
    assign  image_0_835[31:24]   = Image[923];
    assign  image_0_835[23:16]   = Image[953];
    assign  image_0_835[15:8]    = Image[954];
    assign  image_0_835[7:0]     = Image[955];

    assign  image_0_836[71:64]   = Image[890];
    assign  image_0_836[63:56]   = Image[891];
    assign  image_0_836[55:48]   = Image[892];
    assign  image_0_836[47:40]   = Image[922];
    assign  image_0_836[39:32]   = Image[923];
    assign  image_0_836[31:24]   = Image[924];
    assign  image_0_836[23:16]   = Image[954];
    assign  image_0_836[15:8]    = Image[955];
    assign  image_0_836[7:0]     = Image[956];

    assign  image_0_837[71:64]   = Image[891];
    assign  image_0_837[63:56]   = Image[892];
    assign  image_0_837[55:48]   = Image[893];
    assign  image_0_837[47:40]   = Image[923];
    assign  image_0_837[39:32]   = Image[924];
    assign  image_0_837[31:24]   = Image[925];
    assign  image_0_837[23:16]   = Image[955];
    assign  image_0_837[15:8]    = Image[956];
    assign  image_0_837[7:0]     = Image[957];

    assign  image_0_838[71:64]   = Image[892];
    assign  image_0_838[63:56]   = Image[893];
    assign  image_0_838[55:48]   = Image[894];
    assign  image_0_838[47:40]   = Image[924];
    assign  image_0_838[39:32]   = Image[925];
    assign  image_0_838[31:24]   = Image[926];
    assign  image_0_838[23:16]   = Image[956];
    assign  image_0_838[15:8]    = Image[957];
    assign  image_0_838[7:0]     = Image[958];

    assign  image_0_839[71:64]   = Image[893];
    assign  image_0_839[63:56]   = Image[894];
    assign  image_0_839[55:48]   = Image[895];
    assign  image_0_839[47:40]   = Image[925];
    assign  image_0_839[39:32]   = Image[926];
    assign  image_0_839[31:24]   = Image[927];
    assign  image_0_839[23:16]   = Image[957];
    assign  image_0_839[15:8]    = Image[958];
    assign  image_0_839[7:0]     = Image[959];

    assign  image_0_840[71:64]   = Image[896];
    assign  image_0_840[63:56]   = Image[897];
    assign  image_0_840[55:48]   = Image[898];
    assign  image_0_840[47:40]   = Image[928];
    assign  image_0_840[39:32]   = Image[929];
    assign  image_0_840[31:24]   = Image[930];
    assign  image_0_840[23:16]   = Image[960];
    assign  image_0_840[15:8]    = Image[961];
    assign  image_0_840[7:0]     = Image[962];

    assign  image_0_841[71:64]   = Image[897];
    assign  image_0_841[63:56]   = Image[898];
    assign  image_0_841[55:48]   = Image[899];
    assign  image_0_841[47:40]   = Image[929];
    assign  image_0_841[39:32]   = Image[930];
    assign  image_0_841[31:24]   = Image[931];
    assign  image_0_841[23:16]   = Image[961];
    assign  image_0_841[15:8]    = Image[962];
    assign  image_0_841[7:0]     = Image[963];

    assign  image_0_842[71:64]   = Image[898];
    assign  image_0_842[63:56]   = Image[899];
    assign  image_0_842[55:48]   = Image[900];
    assign  image_0_842[47:40]   = Image[930];
    assign  image_0_842[39:32]   = Image[931];
    assign  image_0_842[31:24]   = Image[932];
    assign  image_0_842[23:16]   = Image[962];
    assign  image_0_842[15:8]    = Image[963];
    assign  image_0_842[7:0]     = Image[964];

    assign  image_0_843[71:64]   = Image[899];
    assign  image_0_843[63:56]   = Image[900];
    assign  image_0_843[55:48]   = Image[901];
    assign  image_0_843[47:40]   = Image[931];
    assign  image_0_843[39:32]   = Image[932];
    assign  image_0_843[31:24]   = Image[933];
    assign  image_0_843[23:16]   = Image[963];
    assign  image_0_843[15:8]    = Image[964];
    assign  image_0_843[7:0]     = Image[965];

    assign  image_0_844[71:64]   = Image[900];
    assign  image_0_844[63:56]   = Image[901];
    assign  image_0_844[55:48]   = Image[902];
    assign  image_0_844[47:40]   = Image[932];
    assign  image_0_844[39:32]   = Image[933];
    assign  image_0_844[31:24]   = Image[934];
    assign  image_0_844[23:16]   = Image[964];
    assign  image_0_844[15:8]    = Image[965];
    assign  image_0_844[7:0]     = Image[966];

    assign  image_0_845[71:64]   = Image[901];
    assign  image_0_845[63:56]   = Image[902];
    assign  image_0_845[55:48]   = Image[903];
    assign  image_0_845[47:40]   = Image[933];
    assign  image_0_845[39:32]   = Image[934];
    assign  image_0_845[31:24]   = Image[935];
    assign  image_0_845[23:16]   = Image[965];
    assign  image_0_845[15:8]    = Image[966];
    assign  image_0_845[7:0]     = Image[967];

    assign  image_0_846[71:64]   = Image[902];
    assign  image_0_846[63:56]   = Image[903];
    assign  image_0_846[55:48]   = Image[904];
    assign  image_0_846[47:40]   = Image[934];
    assign  image_0_846[39:32]   = Image[935];
    assign  image_0_846[31:24]   = Image[936];
    assign  image_0_846[23:16]   = Image[966];
    assign  image_0_846[15:8]    = Image[967];
    assign  image_0_846[7:0]     = Image[968];

    assign  image_0_847[71:64]   = Image[903];
    assign  image_0_847[63:56]   = Image[904];
    assign  image_0_847[55:48]   = Image[905];
    assign  image_0_847[47:40]   = Image[935];
    assign  image_0_847[39:32]   = Image[936];
    assign  image_0_847[31:24]   = Image[937];
    assign  image_0_847[23:16]   = Image[967];
    assign  image_0_847[15:8]    = Image[968];
    assign  image_0_847[7:0]     = Image[969];

    assign  image_0_848[71:64]   = Image[904];
    assign  image_0_848[63:56]   = Image[905];
    assign  image_0_848[55:48]   = Image[906];
    assign  image_0_848[47:40]   = Image[936];
    assign  image_0_848[39:32]   = Image[937];
    assign  image_0_848[31:24]   = Image[938];
    assign  image_0_848[23:16]   = Image[968];
    assign  image_0_848[15:8]    = Image[969];
    assign  image_0_848[7:0]     = Image[970];

    assign  image_0_849[71:64]   = Image[905];
    assign  image_0_849[63:56]   = Image[906];
    assign  image_0_849[55:48]   = Image[907];
    assign  image_0_849[47:40]   = Image[937];
    assign  image_0_849[39:32]   = Image[938];
    assign  image_0_849[31:24]   = Image[939];
    assign  image_0_849[23:16]   = Image[969];
    assign  image_0_849[15:8]    = Image[970];
    assign  image_0_849[7:0]     = Image[971];

    assign  image_0_850[71:64]   = Image[906];
    assign  image_0_850[63:56]   = Image[907];
    assign  image_0_850[55:48]   = Image[908];
    assign  image_0_850[47:40]   = Image[938];
    assign  image_0_850[39:32]   = Image[939];
    assign  image_0_850[31:24]   = Image[940];
    assign  image_0_850[23:16]   = Image[970];
    assign  image_0_850[15:8]    = Image[971];
    assign  image_0_850[7:0]     = Image[972];

    assign  image_0_851[71:64]   = Image[907];
    assign  image_0_851[63:56]   = Image[908];
    assign  image_0_851[55:48]   = Image[909];
    assign  image_0_851[47:40]   = Image[939];
    assign  image_0_851[39:32]   = Image[940];
    assign  image_0_851[31:24]   = Image[941];
    assign  image_0_851[23:16]   = Image[971];
    assign  image_0_851[15:8]    = Image[972];
    assign  image_0_851[7:0]     = Image[973];

    assign  image_0_852[71:64]   = Image[908];
    assign  image_0_852[63:56]   = Image[909];
    assign  image_0_852[55:48]   = Image[910];
    assign  image_0_852[47:40]   = Image[940];
    assign  image_0_852[39:32]   = Image[941];
    assign  image_0_852[31:24]   = Image[942];
    assign  image_0_852[23:16]   = Image[972];
    assign  image_0_852[15:8]    = Image[973];
    assign  image_0_852[7:0]     = Image[974];

    assign  image_0_853[71:64]   = Image[909];
    assign  image_0_853[63:56]   = Image[910];
    assign  image_0_853[55:48]   = Image[911];
    assign  image_0_853[47:40]   = Image[941];
    assign  image_0_853[39:32]   = Image[942];
    assign  image_0_853[31:24]   = Image[943];
    assign  image_0_853[23:16]   = Image[973];
    assign  image_0_853[15:8]    = Image[974];
    assign  image_0_853[7:0]     = Image[975];

    assign  image_0_854[71:64]   = Image[910];
    assign  image_0_854[63:56]   = Image[911];
    assign  image_0_854[55:48]   = Image[912];
    assign  image_0_854[47:40]   = Image[942];
    assign  image_0_854[39:32]   = Image[943];
    assign  image_0_854[31:24]   = Image[944];
    assign  image_0_854[23:16]   = Image[974];
    assign  image_0_854[15:8]    = Image[975];
    assign  image_0_854[7:0]     = Image[976];

    assign  image_0_855[71:64]   = Image[911];
    assign  image_0_855[63:56]   = Image[912];
    assign  image_0_855[55:48]   = Image[913];
    assign  image_0_855[47:40]   = Image[943];
    assign  image_0_855[39:32]   = Image[944];
    assign  image_0_855[31:24]   = Image[945];
    assign  image_0_855[23:16]   = Image[975];
    assign  image_0_855[15:8]    = Image[976];
    assign  image_0_855[7:0]     = Image[977];

    assign  image_0_856[71:64]   = Image[912];
    assign  image_0_856[63:56]   = Image[913];
    assign  image_0_856[55:48]   = Image[914];
    assign  image_0_856[47:40]   = Image[944];
    assign  image_0_856[39:32]   = Image[945];
    assign  image_0_856[31:24]   = Image[946];
    assign  image_0_856[23:16]   = Image[976];
    assign  image_0_856[15:8]    = Image[977];
    assign  image_0_856[7:0]     = Image[978];

    assign  image_0_857[71:64]   = Image[913];
    assign  image_0_857[63:56]   = Image[914];
    assign  image_0_857[55:48]   = Image[915];
    assign  image_0_857[47:40]   = Image[945];
    assign  image_0_857[39:32]   = Image[946];
    assign  image_0_857[31:24]   = Image[947];
    assign  image_0_857[23:16]   = Image[977];
    assign  image_0_857[15:8]    = Image[978];
    assign  image_0_857[7:0]     = Image[979];

    assign  image_0_858[71:64]   = Image[914];
    assign  image_0_858[63:56]   = Image[915];
    assign  image_0_858[55:48]   = Image[916];
    assign  image_0_858[47:40]   = Image[946];
    assign  image_0_858[39:32]   = Image[947];
    assign  image_0_858[31:24]   = Image[948];
    assign  image_0_858[23:16]   = Image[978];
    assign  image_0_858[15:8]    = Image[979];
    assign  image_0_858[7:0]     = Image[980];

    assign  image_0_859[71:64]   = Image[915];
    assign  image_0_859[63:56]   = Image[916];
    assign  image_0_859[55:48]   = Image[917];
    assign  image_0_859[47:40]   = Image[947];
    assign  image_0_859[39:32]   = Image[948];
    assign  image_0_859[31:24]   = Image[949];
    assign  image_0_859[23:16]   = Image[979];
    assign  image_0_859[15:8]    = Image[980];
    assign  image_0_859[7:0]     = Image[981];

    assign  image_0_860[71:64]   = Image[916];
    assign  image_0_860[63:56]   = Image[917];
    assign  image_0_860[55:48]   = Image[918];
    assign  image_0_860[47:40]   = Image[948];
    assign  image_0_860[39:32]   = Image[949];
    assign  image_0_860[31:24]   = Image[950];
    assign  image_0_860[23:16]   = Image[980];
    assign  image_0_860[15:8]    = Image[981];
    assign  image_0_860[7:0]     = Image[982];

    assign  image_0_861[71:64]   = Image[917];
    assign  image_0_861[63:56]   = Image[918];
    assign  image_0_861[55:48]   = Image[919];
    assign  image_0_861[47:40]   = Image[949];
    assign  image_0_861[39:32]   = Image[950];
    assign  image_0_861[31:24]   = Image[951];
    assign  image_0_861[23:16]   = Image[981];
    assign  image_0_861[15:8]    = Image[982];
    assign  image_0_861[7:0]     = Image[983];

    assign  image_0_862[71:64]   = Image[918];
    assign  image_0_862[63:56]   = Image[919];
    assign  image_0_862[55:48]   = Image[920];
    assign  image_0_862[47:40]   = Image[950];
    assign  image_0_862[39:32]   = Image[951];
    assign  image_0_862[31:24]   = Image[952];
    assign  image_0_862[23:16]   = Image[982];
    assign  image_0_862[15:8]    = Image[983];
    assign  image_0_862[7:0]     = Image[984];

    assign  image_0_863[71:64]   = Image[919];
    assign  image_0_863[63:56]   = Image[920];
    assign  image_0_863[55:48]   = Image[921];
    assign  image_0_863[47:40]   = Image[951];
    assign  image_0_863[39:32]   = Image[952];
    assign  image_0_863[31:24]   = Image[953];
    assign  image_0_863[23:16]   = Image[983];
    assign  image_0_863[15:8]    = Image[984];
    assign  image_0_863[7:0]     = Image[985];

    assign  image_0_864[71:64]   = Image[920];
    assign  image_0_864[63:56]   = Image[921];
    assign  image_0_864[55:48]   = Image[922];
    assign  image_0_864[47:40]   = Image[952];
    assign  image_0_864[39:32]   = Image[953];
    assign  image_0_864[31:24]   = Image[954];
    assign  image_0_864[23:16]   = Image[984];
    assign  image_0_864[15:8]    = Image[985];
    assign  image_0_864[7:0]     = Image[986];

    assign  image_0_865[71:64]   = Image[921];
    assign  image_0_865[63:56]   = Image[922];
    assign  image_0_865[55:48]   = Image[923];
    assign  image_0_865[47:40]   = Image[953];
    assign  image_0_865[39:32]   = Image[954];
    assign  image_0_865[31:24]   = Image[955];
    assign  image_0_865[23:16]   = Image[985];
    assign  image_0_865[15:8]    = Image[986];
    assign  image_0_865[7:0]     = Image[987];

    assign  image_0_866[71:64]   = Image[922];
    assign  image_0_866[63:56]   = Image[923];
    assign  image_0_866[55:48]   = Image[924];
    assign  image_0_866[47:40]   = Image[954];
    assign  image_0_866[39:32]   = Image[955];
    assign  image_0_866[31:24]   = Image[956];
    assign  image_0_866[23:16]   = Image[986];
    assign  image_0_866[15:8]    = Image[987];
    assign  image_0_866[7:0]     = Image[988];

    assign  image_0_867[71:64]   = Image[923];
    assign  image_0_867[63:56]   = Image[924];
    assign  image_0_867[55:48]   = Image[925];
    assign  image_0_867[47:40]   = Image[955];
    assign  image_0_867[39:32]   = Image[956];
    assign  image_0_867[31:24]   = Image[957];
    assign  image_0_867[23:16]   = Image[987];
    assign  image_0_867[15:8]    = Image[988];
    assign  image_0_867[7:0]     = Image[989];

    assign  image_0_868[71:64]   = Image[924];
    assign  image_0_868[63:56]   = Image[925];
    assign  image_0_868[55:48]   = Image[926];
    assign  image_0_868[47:40]   = Image[956];
    assign  image_0_868[39:32]   = Image[957];
    assign  image_0_868[31:24]   = Image[958];
    assign  image_0_868[23:16]   = Image[988];
    assign  image_0_868[15:8]    = Image[989];
    assign  image_0_868[7:0]     = Image[990];

    assign  image_0_869[71:64]   = Image[925];
    assign  image_0_869[63:56]   = Image[926];
    assign  image_0_869[55:48]   = Image[927];
    assign  image_0_869[47:40]   = Image[957];
    assign  image_0_869[39:32]   = Image[958];
    assign  image_0_869[31:24]   = Image[959];
    assign  image_0_869[23:16]   = Image[989];
    assign  image_0_869[15:8]    = Image[990];
    assign  image_0_869[7:0]     = Image[991];

    assign  image_0_870[71:64]   = Image[928];
    assign  image_0_870[63:56]   = Image[929];
    assign  image_0_870[55:48]   = Image[930];
    assign  image_0_870[47:40]   = Image[960];
    assign  image_0_870[39:32]   = Image[961];
    assign  image_0_870[31:24]   = Image[962];
    assign  image_0_870[23:16]   = Image[992];
    assign  image_0_870[15:8]    = Image[993];
    assign  image_0_870[7:0]     = Image[994];

    assign  image_0_871[71:64]   = Image[929];
    assign  image_0_871[63:56]   = Image[930];
    assign  image_0_871[55:48]   = Image[931];
    assign  image_0_871[47:40]   = Image[961];
    assign  image_0_871[39:32]   = Image[962];
    assign  image_0_871[31:24]   = Image[963];
    assign  image_0_871[23:16]   = Image[993];
    assign  image_0_871[15:8]    = Image[994];
    assign  image_0_871[7:0]     = Image[995];

    assign  image_0_872[71:64]   = Image[930];
    assign  image_0_872[63:56]   = Image[931];
    assign  image_0_872[55:48]   = Image[932];
    assign  image_0_872[47:40]   = Image[962];
    assign  image_0_872[39:32]   = Image[963];
    assign  image_0_872[31:24]   = Image[964];
    assign  image_0_872[23:16]   = Image[994];
    assign  image_0_872[15:8]    = Image[995];
    assign  image_0_872[7:0]     = Image[996];

    assign  image_0_873[71:64]   = Image[931];
    assign  image_0_873[63:56]   = Image[932];
    assign  image_0_873[55:48]   = Image[933];
    assign  image_0_873[47:40]   = Image[963];
    assign  image_0_873[39:32]   = Image[964];
    assign  image_0_873[31:24]   = Image[965];
    assign  image_0_873[23:16]   = Image[995];
    assign  image_0_873[15:8]    = Image[996];
    assign  image_0_873[7:0]     = Image[997];

    assign  image_0_874[71:64]   = Image[932];
    assign  image_0_874[63:56]   = Image[933];
    assign  image_0_874[55:48]   = Image[934];
    assign  image_0_874[47:40]   = Image[964];
    assign  image_0_874[39:32]   = Image[965];
    assign  image_0_874[31:24]   = Image[966];
    assign  image_0_874[23:16]   = Image[996];
    assign  image_0_874[15:8]    = Image[997];
    assign  image_0_874[7:0]     = Image[998];

    assign  image_0_875[71:64]   = Image[933];
    assign  image_0_875[63:56]   = Image[934];
    assign  image_0_875[55:48]   = Image[935];
    assign  image_0_875[47:40]   = Image[965];
    assign  image_0_875[39:32]   = Image[966];
    assign  image_0_875[31:24]   = Image[967];
    assign  image_0_875[23:16]   = Image[997];
    assign  image_0_875[15:8]    = Image[998];
    assign  image_0_875[7:0]     = Image[999];

    assign  image_0_876[71:64]   = Image[934];
    assign  image_0_876[63:56]   = Image[935];
    assign  image_0_876[55:48]   = Image[936];
    assign  image_0_876[47:40]   = Image[966];
    assign  image_0_876[39:32]   = Image[967];
    assign  image_0_876[31:24]   = Image[968];
    assign  image_0_876[23:16]   = Image[998];
    assign  image_0_876[15:8]    = Image[999];
    assign  image_0_876[7:0]     = Image[1000];

    assign  image_0_877[71:64]   = Image[935];
    assign  image_0_877[63:56]   = Image[936];
    assign  image_0_877[55:48]   = Image[937];
    assign  image_0_877[47:40]   = Image[967];
    assign  image_0_877[39:32]   = Image[968];
    assign  image_0_877[31:24]   = Image[969];
    assign  image_0_877[23:16]   = Image[999];
    assign  image_0_877[15:8]    = Image[1000];
    assign  image_0_877[7:0]     = Image[1001];

    assign  image_0_878[71:64]   = Image[936];
    assign  image_0_878[63:56]   = Image[937];
    assign  image_0_878[55:48]   = Image[938];
    assign  image_0_878[47:40]   = Image[968];
    assign  image_0_878[39:32]   = Image[969];
    assign  image_0_878[31:24]   = Image[970];
    assign  image_0_878[23:16]   = Image[1000];
    assign  image_0_878[15:8]    = Image[1001];
    assign  image_0_878[7:0]     = Image[1002];

    assign  image_0_879[71:64]   = Image[937];
    assign  image_0_879[63:56]   = Image[938];
    assign  image_0_879[55:48]   = Image[939];
    assign  image_0_879[47:40]   = Image[969];
    assign  image_0_879[39:32]   = Image[970];
    assign  image_0_879[31:24]   = Image[971];
    assign  image_0_879[23:16]   = Image[1001];
    assign  image_0_879[15:8]    = Image[1002];
    assign  image_0_879[7:0]     = Image[1003];

    assign  image_0_880[71:64]   = Image[938];
    assign  image_0_880[63:56]   = Image[939];
    assign  image_0_880[55:48]   = Image[940];
    assign  image_0_880[47:40]   = Image[970];
    assign  image_0_880[39:32]   = Image[971];
    assign  image_0_880[31:24]   = Image[972];
    assign  image_0_880[23:16]   = Image[1002];
    assign  image_0_880[15:8]    = Image[1003];
    assign  image_0_880[7:0]     = Image[1004];

    assign  image_0_881[71:64]   = Image[939];
    assign  image_0_881[63:56]   = Image[940];
    assign  image_0_881[55:48]   = Image[941];
    assign  image_0_881[47:40]   = Image[971];
    assign  image_0_881[39:32]   = Image[972];
    assign  image_0_881[31:24]   = Image[973];
    assign  image_0_881[23:16]   = Image[1003];
    assign  image_0_881[15:8]    = Image[1004];
    assign  image_0_881[7:0]     = Image[1005];

    assign  image_0_882[71:64]   = Image[940];
    assign  image_0_882[63:56]   = Image[941];
    assign  image_0_882[55:48]   = Image[942];
    assign  image_0_882[47:40]   = Image[972];
    assign  image_0_882[39:32]   = Image[973];
    assign  image_0_882[31:24]   = Image[974];
    assign  image_0_882[23:16]   = Image[1004];
    assign  image_0_882[15:8]    = Image[1005];
    assign  image_0_882[7:0]     = Image[1006];

    assign  image_0_883[71:64]   = Image[941];
    assign  image_0_883[63:56]   = Image[942];
    assign  image_0_883[55:48]   = Image[943];
    assign  image_0_883[47:40]   = Image[973];
    assign  image_0_883[39:32]   = Image[974];
    assign  image_0_883[31:24]   = Image[975];
    assign  image_0_883[23:16]   = Image[1005];
    assign  image_0_883[15:8]    = Image[1006];
    assign  image_0_883[7:0]     = Image[1007];

    assign  image_0_884[71:64]   = Image[942];
    assign  image_0_884[63:56]   = Image[943];
    assign  image_0_884[55:48]   = Image[944];
    assign  image_0_884[47:40]   = Image[974];
    assign  image_0_884[39:32]   = Image[975];
    assign  image_0_884[31:24]   = Image[976];
    assign  image_0_884[23:16]   = Image[1006];
    assign  image_0_884[15:8]    = Image[1007];
    assign  image_0_884[7:0]     = Image[1008];

    assign  image_0_885[71:64]   = Image[943];
    assign  image_0_885[63:56]   = Image[944];
    assign  image_0_885[55:48]   = Image[945];
    assign  image_0_885[47:40]   = Image[975];
    assign  image_0_885[39:32]   = Image[976];
    assign  image_0_885[31:24]   = Image[977];
    assign  image_0_885[23:16]   = Image[1007];
    assign  image_0_885[15:8]    = Image[1008];
    assign  image_0_885[7:0]     = Image[1009];

    assign  image_0_886[71:64]   = Image[944];
    assign  image_0_886[63:56]   = Image[945];
    assign  image_0_886[55:48]   = Image[946];
    assign  image_0_886[47:40]   = Image[976];
    assign  image_0_886[39:32]   = Image[977];
    assign  image_0_886[31:24]   = Image[978];
    assign  image_0_886[23:16]   = Image[1008];
    assign  image_0_886[15:8]    = Image[1009];
    assign  image_0_886[7:0]     = Image[1010];

    assign  image_0_887[71:64]   = Image[945];
    assign  image_0_887[63:56]   = Image[946];
    assign  image_0_887[55:48]   = Image[947];
    assign  image_0_887[47:40]   = Image[977];
    assign  image_0_887[39:32]   = Image[978];
    assign  image_0_887[31:24]   = Image[979];
    assign  image_0_887[23:16]   = Image[1009];
    assign  image_0_887[15:8]    = Image[1010];
    assign  image_0_887[7:0]     = Image[1011];

    assign  image_0_888[71:64]   = Image[946];
    assign  image_0_888[63:56]   = Image[947];
    assign  image_0_888[55:48]   = Image[948];
    assign  image_0_888[47:40]   = Image[978];
    assign  image_0_888[39:32]   = Image[979];
    assign  image_0_888[31:24]   = Image[980];
    assign  image_0_888[23:16]   = Image[1010];
    assign  image_0_888[15:8]    = Image[1011];
    assign  image_0_888[7:0]     = Image[1012];

    assign  image_0_889[71:64]   = Image[947];
    assign  image_0_889[63:56]   = Image[948];
    assign  image_0_889[55:48]   = Image[949];
    assign  image_0_889[47:40]   = Image[979];
    assign  image_0_889[39:32]   = Image[980];
    assign  image_0_889[31:24]   = Image[981];
    assign  image_0_889[23:16]   = Image[1011];
    assign  image_0_889[15:8]    = Image[1012];
    assign  image_0_889[7:0]     = Image[1013];

    assign  image_0_890[71:64]   = Image[948];
    assign  image_0_890[63:56]   = Image[949];
    assign  image_0_890[55:48]   = Image[950];
    assign  image_0_890[47:40]   = Image[980];
    assign  image_0_890[39:32]   = Image[981];
    assign  image_0_890[31:24]   = Image[982];
    assign  image_0_890[23:16]   = Image[1012];
    assign  image_0_890[15:8]    = Image[1013];
    assign  image_0_890[7:0]     = Image[1014];

    assign  image_0_891[71:64]   = Image[949];
    assign  image_0_891[63:56]   = Image[950];
    assign  image_0_891[55:48]   = Image[951];
    assign  image_0_891[47:40]   = Image[981];
    assign  image_0_891[39:32]   = Image[982];
    assign  image_0_891[31:24]   = Image[983];
    assign  image_0_891[23:16]   = Image[1013];
    assign  image_0_891[15:8]    = Image[1014];
    assign  image_0_891[7:0]     = Image[1015];

    assign  image_0_892[71:64]   = Image[950];
    assign  image_0_892[63:56]   = Image[951];
    assign  image_0_892[55:48]   = Image[952];
    assign  image_0_892[47:40]   = Image[982];
    assign  image_0_892[39:32]   = Image[983];
    assign  image_0_892[31:24]   = Image[984];
    assign  image_0_892[23:16]   = Image[1014];
    assign  image_0_892[15:8]    = Image[1015];
    assign  image_0_892[7:0]     = Image[1016];

    assign  image_0_893[71:64]   = Image[951];
    assign  image_0_893[63:56]   = Image[952];
    assign  image_0_893[55:48]   = Image[953];
    assign  image_0_893[47:40]   = Image[983];
    assign  image_0_893[39:32]   = Image[984];
    assign  image_0_893[31:24]   = Image[985];
    assign  image_0_893[23:16]   = Image[1015];
    assign  image_0_893[15:8]    = Image[1016];
    assign  image_0_893[7:0]     = Image[1017];

    assign  image_0_894[71:64]   = Image[952];
    assign  image_0_894[63:56]   = Image[953];
    assign  image_0_894[55:48]   = Image[954];
    assign  image_0_894[47:40]   = Image[984];
    assign  image_0_894[39:32]   = Image[985];
    assign  image_0_894[31:24]   = Image[986];
    assign  image_0_894[23:16]   = Image[1016];
    assign  image_0_894[15:8]    = Image[1017];
    assign  image_0_894[7:0]     = Image[1018];

    assign  image_0_895[71:64]   = Image[953];
    assign  image_0_895[63:56]   = Image[954];
    assign  image_0_895[55:48]   = Image[955];
    assign  image_0_895[47:40]   = Image[985];
    assign  image_0_895[39:32]   = Image[986];
    assign  image_0_895[31:24]   = Image[987];
    assign  image_0_895[23:16]   = Image[1017];
    assign  image_0_895[15:8]    = Image[1018];
    assign  image_0_895[7:0]     = Image[1019];

    assign  image_0_896[71:64]   = Image[954];
    assign  image_0_896[63:56]   = Image[955];
    assign  image_0_896[55:48]   = Image[956];
    assign  image_0_896[47:40]   = Image[986];
    assign  image_0_896[39:32]   = Image[987];
    assign  image_0_896[31:24]   = Image[988];
    assign  image_0_896[23:16]   = Image[1018];
    assign  image_0_896[15:8]    = Image[1019];
    assign  image_0_896[7:0]     = Image[1020];

    assign  image_0_897[71:64]   = Image[955];
    assign  image_0_897[63:56]   = Image[956];
    assign  image_0_897[55:48]   = Image[957];
    assign  image_0_897[47:40]   = Image[987];
    assign  image_0_897[39:32]   = Image[988];
    assign  image_0_897[31:24]   = Image[989];
    assign  image_0_897[23:16]   = Image[1019];
    assign  image_0_897[15:8]    = Image[1020];
    assign  image_0_897[7:0]     = Image[1021];

    assign  image_0_898[71:64]   = Image[956];
    assign  image_0_898[63:56]   = Image[957];
    assign  image_0_898[55:48]   = Image[958];
    assign  image_0_898[47:40]   = Image[988];
    assign  image_0_898[39:32]   = Image[989];
    assign  image_0_898[31:24]   = Image[990];
    assign  image_0_898[23:16]   = Image[1020];
    assign  image_0_898[15:8]    = Image[1021];
    assign  image_0_898[7:0]     = Image[1022];

    assign  image_0_899[71:64]   = Image[957];
    assign  image_0_899[63:56]   = Image[958];
    assign  image_0_899[55:48]   = Image[959];
    assign  image_0_899[47:40]   = Image[989];
    assign  image_0_899[39:32]   = Image[990];
    assign  image_0_899[31:24]   = Image[991];
    assign  image_0_899[23:16]   = Image[1021];
    assign  image_0_899[15:8]    = Image[1022];
    assign  image_0_899[7:0]     = Image[1023];


    assign  filter = Filter; 
    assign  filter_0 = Filter_0;
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////  
wire    [143:0]  image_1_0, image_1_1, image_1_2, image_1_3, image_1_4, image_1_5, image_1_6, image_1_7, image_1_8, image_1_9, image_1_10, image_1_11, image_1_12, image_1_13;
wire    [143:0]  image_1_14, image_1_15, image_1_16, image_1_17, image_1_18, image_1_19, image_1_20, image_1_21, image_1_22, image_1_23, image_1_24, image_1_25, image_1_26, image_1_27;
wire    [143:0]  image_1_28, image_1_29, image_1_30, image_1_31, image_1_32, image_1_33, image_1_34, image_1_35, image_1_36, image_1_37, image_1_38, image_1_39, image_1_40, image_1_41;
wire    [143:0]  image_1_42, image_1_43, image_1_44, image_1_45, image_1_46, image_1_47, image_1_48, image_1_49, image_1_50, image_1_51, image_1_52, image_1_53, image_1_54, image_1_55;
wire    [143:0]  image_1_56, image_1_57, image_1_58, image_1_59, image_1_60, image_1_61, image_1_62, image_1_63, image_1_64, image_1_65, image_1_66, image_1_67, image_1_68, image_1_69;
wire    [143:0]  image_1_70, image_1_71, image_1_72, image_1_73, image_1_74, image_1_75, image_1_76, image_1_77, image_1_78, image_1_79, image_1_80, image_1_81, image_1_82, image_1_83;
wire    [143:0]  image_1_84, image_1_85, image_1_86, image_1_87, image_1_88, image_1_89, image_1_90, image_1_91, image_1_92, image_1_93, image_1_94, image_1_95, image_1_96, image_1_97;
wire    [143:0]  image_1_98, image_1_99, image_1_100, image_1_101, image_1_102, image_1_103, image_1_104, image_1_105, image_1_106, image_1_107, image_1_108, image_1_109, image_1_110, image_1_111;
wire    [143:0]  image_1_112, image_1_113, image_1_114, image_1_115, image_1_116, image_1_117, image_1_118, image_1_119, image_1_120, image_1_121, image_1_122, image_1_123, image_1_124, image_1_125;
wire    [143:0]  image_1_126, image_1_127, image_1_128, image_1_129, image_1_130, image_1_131, image_1_132, image_1_133, image_1_134, image_1_135, image_1_136, image_1_137, image_1_138, image_1_139;
wire    [143:0]  image_1_140, image_1_141, image_1_142, image_1_143, image_1_144, image_1_145, image_1_146, image_1_147, image_1_148, image_1_149, image_1_150, image_1_151, image_1_152, image_1_153;
wire    [143:0]  image_1_154, image_1_155, image_1_156, image_1_157, image_1_158, image_1_159, image_1_160, image_1_161, image_1_162, image_1_163, image_1_164, image_1_165, image_1_166, image_1_167;
wire    [143:0]  image_1_168, image_1_169, image_1_170, image_1_171, image_1_172, image_1_173, image_1_174, image_1_175, image_1_176, image_1_177, image_1_178, image_1_179, image_1_180, image_1_181;
wire    [143:0]  image_1_182, image_1_183, image_1_184, image_1_185, image_1_186, image_1_187, image_1_188, image_1_189, image_1_190, image_1_191, image_1_192, image_1_193, image_1_194, image_1_195;
wire    [143:0]  image_1_196, image_1_197, image_1_198, image_1_199, image_1_200, image_1_201, image_1_202, image_1_203, image_1_204, image_1_205, image_1_206, image_1_207, image_1_208, image_1_209;
wire    [143:0]  image_1_210, image_1_211, image_1_212, image_1_213, image_1_214, image_1_215, image_1_216, image_1_217, image_1_218, image_1_219, image_1_220, image_1_221, image_1_222, image_1_223;
wire    [143:0]  image_1_224, image_1_225, image_1_226, image_1_227, image_1_228, image_1_229, image_1_230, image_1_231, image_1_232, image_1_233, image_1_234, image_1_235, image_1_236, image_1_237;
wire    [143:0]  image_1_238, image_1_239, image_1_240, image_1_241, image_1_242, image_1_243, image_1_244, image_1_245, image_1_246, image_1_247, image_1_248, image_1_249, image_1_250, image_1_251;
wire    [143:0]  image_1_252, image_1_253, image_1_254, image_1_255, image_1_256, image_1_257, image_1_258, image_1_259, image_1_260, image_1_261, image_1_262, image_1_263, image_1_264, image_1_265;
wire    [143:0]  image_1_266, image_1_267, image_1_268, image_1_269, image_1_270, image_1_271, image_1_272, image_1_273, image_1_274, image_1_275, image_1_276, image_1_277, image_1_278, image_1_279;
wire    [143:0]  image_1_280, image_1_281, image_1_282, image_1_283, image_1_284, image_1_285, image_1_286, image_1_287, image_1_288, image_1_289, image_1_290, image_1_291, image_1_292, image_1_293;
wire    [143:0]  image_1_294, image_1_295, image_1_296, image_1_297, image_1_298, image_1_299, image_1_300, image_1_301, image_1_302, image_1_303, image_1_304, image_1_305, image_1_306, image_1_307;
wire    [143:0]  image_1_308, image_1_309, image_1_310, image_1_311, image_1_312, image_1_313, image_1_314, image_1_315, image_1_316, image_1_317, image_1_318, image_1_319, image_1_320, image_1_321;
wire    [143:0]  image_1_322, image_1_323, image_1_324, image_1_325, image_1_326, image_1_327, image_1_328, image_1_329, image_1_330, image_1_331, image_1_332, image_1_333, image_1_334, image_1_335;
wire    [143:0]  image_1_336, image_1_337, image_1_338, image_1_339, image_1_340, image_1_341, image_1_342, image_1_343, image_1_344, image_1_345, image_1_346, image_1_347, image_1_348, image_1_349;
wire    [143:0]  image_1_350, image_1_351, image_1_352, image_1_353, image_1_354, image_1_355, image_1_356, image_1_357, image_1_358, image_1_359, image_1_360, image_1_361, image_1_362, image_1_363;
wire    [143:0]  image_1_364, image_1_365, image_1_366, image_1_367, image_1_368, image_1_369, image_1_370, image_1_371, image_1_372, image_1_373, image_1_374, image_1_375, image_1_376, image_1_377;
wire    [143:0]  image_1_378, image_1_379, image_1_380, image_1_381, image_1_382, image_1_383, image_1_384, image_1_385, image_1_386, image_1_387, image_1_388, image_1_389, image_1_390, image_1_391;
wire    [143:0]  image_1_392, image_1_393, image_1_394, image_1_395, image_1_396, image_1_397, image_1_398, image_1_399, image_1_400, image_1_401, image_1_402, image_1_403, image_1_404, image_1_405;
wire    [143:0]  image_1_406, image_1_407, image_1_408, image_1_409, image_1_410, image_1_411, image_1_412, image_1_413, image_1_414, image_1_415, image_1_416, image_1_417, image_1_418, image_1_419;
wire    [143:0]  image_1_420, image_1_421, image_1_422, image_1_423, image_1_424, image_1_425, image_1_426, image_1_427, image_1_428, image_1_429, image_1_430, image_1_431, image_1_432, image_1_433;
wire    [143:0]  image_1_434, image_1_435, image_1_436, image_1_437, image_1_438, image_1_439, image_1_440, image_1_441, image_1_442, image_1_443, image_1_444, image_1_445, image_1_446, image_1_447;
wire    [143:0]  image_1_448, image_1_449, image_1_450, image_1_451, image_1_452, image_1_453, image_1_454, image_1_455, image_1_456, image_1_457, image_1_458, image_1_459, image_1_460, image_1_461;
wire    [143:0]  image_1_462, image_1_463, image_1_464, image_1_465, image_1_466, image_1_467, image_1_468, image_1_469, image_1_470, image_1_471, image_1_472, image_1_473, image_1_474, image_1_475;
wire    [143:0]  image_1_476, image_1_477, image_1_478, image_1_479, image_1_480, image_1_481, image_1_482, image_1_483, image_1_484, image_1_485, image_1_486, image_1_487, image_1_488, image_1_489;
wire    [143:0]  image_1_490, image_1_491, image_1_492, image_1_493, image_1_494, image_1_495, image_1_496, image_1_497, image_1_498, image_1_499, image_1_500, image_1_501, image_1_502, image_1_503;
wire    [143:0]  image_1_504, image_1_505, image_1_506, image_1_507, image_1_508, image_1_509, image_1_510, image_1_511, image_1_512, image_1_513, image_1_514, image_1_515, image_1_516, image_1_517;
wire    [143:0]  image_1_518, image_1_519, image_1_520, image_1_521, image_1_522, image_1_523, image_1_524, image_1_525, image_1_526, image_1_527, image_1_528, image_1_529, image_1_530, image_1_531;
wire    [143:0]  image_1_532, image_1_533, image_1_534, image_1_535, image_1_536, image_1_537, image_1_538, image_1_539, image_1_540, image_1_541, image_1_542, image_1_543, image_1_544, image_1_545;
wire    [143:0]  image_1_546, image_1_547, image_1_548, image_1_549, image_1_550, image_1_551, image_1_552, image_1_553, image_1_554, image_1_555, image_1_556, image_1_557, image_1_558, image_1_559;
wire    [143:0]  image_1_560, image_1_561, image_1_562, image_1_563, image_1_564, image_1_565, image_1_566, image_1_567, image_1_568, image_1_569, image_1_570, image_1_571, image_1_572, image_1_573;
wire    [143:0]  image_1_574, image_1_575, image_1_576, image_1_577, image_1_578, image_1_579, image_1_580, image_1_581, image_1_582, image_1_583, image_1_584, image_1_585, image_1_586, image_1_587;
wire    [143:0]  image_1_588, image_1_589, image_1_590, image_1_591, image_1_592, image_1_593, image_1_594, image_1_595, image_1_596, image_1_597, image_1_598, image_1_599, image_1_600, image_1_601;
wire    [143:0]  image_1_602, image_1_603, image_1_604, image_1_605, image_1_606, image_1_607, image_1_608, image_1_609, image_1_610, image_1_611, image_1_612, image_1_613, image_1_614, image_1_615;
wire    [143:0]  image_1_616, image_1_617, image_1_618, image_1_619, image_1_620, image_1_621, image_1_622, image_1_623, image_1_624, image_1_625, image_1_626, image_1_627, image_1_628, image_1_629;
wire    [143:0]  image_1_630, image_1_631, image_1_632, image_1_633, image_1_634, image_1_635, image_1_636, image_1_637, image_1_638, image_1_639, image_1_640, image_1_641, image_1_642, image_1_643;
wire    [143:0]  image_1_644, image_1_645, image_1_646, image_1_647, image_1_648, image_1_649, image_1_650, image_1_651, image_1_652, image_1_653, image_1_654, image_1_655, image_1_656, image_1_657;
wire    [143:0]  image_1_658, image_1_659, image_1_660, image_1_661, image_1_662, image_1_663, image_1_664, image_1_665, image_1_666, image_1_667, image_1_668, image_1_669, image_1_670, image_1_671;
wire    [143:0]  image_1_672, image_1_673, image_1_674, image_1_675, image_1_676, image_1_677, image_1_678, image_1_679, image_1_680, image_1_681, image_1_682, image_1_683, image_1_684, image_1_685;
wire    [143:0]  image_1_686, image_1_687, image_1_688, image_1_689, image_1_690, image_1_691, image_1_692, image_1_693, image_1_694, image_1_695, image_1_696, image_1_697, image_1_698, image_1_699;
wire    [143:0]  image_1_700, image_1_701, image_1_702, image_1_703, image_1_704, image_1_705, image_1_706, image_1_707, image_1_708, image_1_709, image_1_710, image_1_711, image_1_712, image_1_713;
wire    [143:0]  image_1_714, image_1_715, image_1_716, image_1_717, image_1_718, image_1_719, image_1_720, image_1_721, image_1_722, image_1_723, image_1_724, image_1_725, image_1_726, image_1_727;
wire    [143:0]  image_1_728, image_1_729, image_1_730, image_1_731, image_1_732, image_1_733, image_1_734, image_1_735, image_1_736, image_1_737, image_1_738, image_1_739, image_1_740, image_1_741;
wire    [143:0]  image_1_742, image_1_743, image_1_744, image_1_745, image_1_746, image_1_747, image_1_748, image_1_749, image_1_750, image_1_751, image_1_752, image_1_753, image_1_754, image_1_755;
wire    [143:0]  image_1_756, image_1_757, image_1_758, image_1_759, image_1_760, image_1_761, image_1_762, image_1_763, image_1_764, image_1_765, image_1_766, image_1_767, image_1_768, image_1_769;
wire    [143:0]  image_1_770, image_1_771, image_1_772, image_1_773, image_1_774, image_1_775, image_1_776, image_1_777, image_1_778, image_1_779, image_1_780, image_1_781, image_1_782, image_1_783;

wire    [31:0]  conv_out_1_0, conv_out_1_1, conv_out_1_2, conv_out_1_3, conv_out_1_4, conv_out_1_5, conv_out_1_6, conv_out_1_7, conv_out_1_8, conv_out_1_9, conv_out_1_10, conv_out_1_11, conv_out_1_12, conv_out_1_13;
wire    [31:0]  conv_out_1_14, conv_out_1_15, conv_out_1_16, conv_out_1_17, conv_out_1_18, conv_out_1_19, conv_out_1_20, conv_out_1_21, conv_out_1_22, conv_out_1_23, conv_out_1_24, conv_out_1_25, conv_out_1_26, conv_out_1_27;
wire    [31:0]  conv_out_1_28, conv_out_1_29, conv_out_1_30, conv_out_1_31, conv_out_1_32, conv_out_1_33, conv_out_1_34, conv_out_1_35, conv_out_1_36, conv_out_1_37, conv_out_1_38, conv_out_1_39, conv_out_1_40, conv_out_1_41;
wire    [31:0]  conv_out_1_42, conv_out_1_43, conv_out_1_44, conv_out_1_45, conv_out_1_46, conv_out_1_47, conv_out_1_48, conv_out_1_49, conv_out_1_50, conv_out_1_51, conv_out_1_52, conv_out_1_53, conv_out_1_54, conv_out_1_55;
wire    [31:0]  conv_out_1_56, conv_out_1_57, conv_out_1_58, conv_out_1_59, conv_out_1_60, conv_out_1_61, conv_out_1_62, conv_out_1_63, conv_out_1_64, conv_out_1_65, conv_out_1_66, conv_out_1_67, conv_out_1_68, conv_out_1_69;
wire    [31:0]  conv_out_1_70, conv_out_1_71, conv_out_1_72, conv_out_1_73, conv_out_1_74, conv_out_1_75, conv_out_1_76, conv_out_1_77, conv_out_1_78, conv_out_1_79, conv_out_1_80, conv_out_1_81, conv_out_1_82, conv_out_1_83;
wire    [31:0]  conv_out_1_84, conv_out_1_85, conv_out_1_86, conv_out_1_87, conv_out_1_88, conv_out_1_89, conv_out_1_90, conv_out_1_91, conv_out_1_92, conv_out_1_93, conv_out_1_94, conv_out_1_95, conv_out_1_96, conv_out_1_97;
wire    [31:0]  conv_out_1_98, conv_out_1_99, conv_out_1_100, conv_out_1_101, conv_out_1_102, conv_out_1_103, conv_out_1_104, conv_out_1_105, conv_out_1_106, conv_out_1_107, conv_out_1_108, conv_out_1_109, conv_out_1_110, conv_out_1_111;
wire    [31:0]  conv_out_1_112, conv_out_1_113, conv_out_1_114, conv_out_1_115, conv_out_1_116, conv_out_1_117, conv_out_1_118, conv_out_1_119, conv_out_1_120, conv_out_1_121, conv_out_1_122, conv_out_1_123, conv_out_1_124, conv_out_1_125;
wire    [31:0]  conv_out_1_126, conv_out_1_127, conv_out_1_128, conv_out_1_129, conv_out_1_130, conv_out_1_131, conv_out_1_132, conv_out_1_133, conv_out_1_134, conv_out_1_135, conv_out_1_136, conv_out_1_137, conv_out_1_138, conv_out_1_139;
wire    [31:0]  conv_out_1_140, conv_out_1_141, conv_out_1_142, conv_out_1_143, conv_out_1_144, conv_out_1_145, conv_out_1_146, conv_out_1_147, conv_out_1_148, conv_out_1_149, conv_out_1_150, conv_out_1_151, conv_out_1_152, conv_out_1_153;
wire    [31:0]  conv_out_1_154, conv_out_1_155, conv_out_1_156, conv_out_1_157, conv_out_1_158, conv_out_1_159, conv_out_1_160, conv_out_1_161, conv_out_1_162, conv_out_1_163, conv_out_1_164, conv_out_1_165, conv_out_1_166, conv_out_1_167;
wire    [31:0]  conv_out_1_168, conv_out_1_169, conv_out_1_170, conv_out_1_171, conv_out_1_172, conv_out_1_173, conv_out_1_174, conv_out_1_175, conv_out_1_176, conv_out_1_177, conv_out_1_178, conv_out_1_179, conv_out_1_180, conv_out_1_181;
wire    [31:0]  conv_out_1_182, conv_out_1_183, conv_out_1_184, conv_out_1_185, conv_out_1_186, conv_out_1_187, conv_out_1_188, conv_out_1_189, conv_out_1_190, conv_out_1_191, conv_out_1_192, conv_out_1_193, conv_out_1_194, conv_out_1_195;
wire    [31:0]  conv_out_1_196, conv_out_1_197, conv_out_1_198, conv_out_1_199, conv_out_1_200, conv_out_1_201, conv_out_1_202, conv_out_1_203, conv_out_1_204, conv_out_1_205, conv_out_1_206, conv_out_1_207, conv_out_1_208, conv_out_1_209;
wire    [31:0]  conv_out_1_210, conv_out_1_211, conv_out_1_212, conv_out_1_213, conv_out_1_214, conv_out_1_215, conv_out_1_216, conv_out_1_217, conv_out_1_218, conv_out_1_219, conv_out_1_220, conv_out_1_221, conv_out_1_222, conv_out_1_223;
wire    [31:0]  conv_out_1_224, conv_out_1_225, conv_out_1_226, conv_out_1_227, conv_out_1_228, conv_out_1_229, conv_out_1_230, conv_out_1_231, conv_out_1_232, conv_out_1_233, conv_out_1_234, conv_out_1_235, conv_out_1_236, conv_out_1_237;
wire    [31:0]  conv_out_1_238, conv_out_1_239, conv_out_1_240, conv_out_1_241, conv_out_1_242, conv_out_1_243, conv_out_1_244, conv_out_1_245, conv_out_1_246, conv_out_1_247, conv_out_1_248, conv_out_1_249, conv_out_1_250, conv_out_1_251;
wire    [31:0]  conv_out_1_252, conv_out_1_253, conv_out_1_254, conv_out_1_255, conv_out_1_256, conv_out_1_257, conv_out_1_258, conv_out_1_259, conv_out_1_260, conv_out_1_261, conv_out_1_262, conv_out_1_263, conv_out_1_264, conv_out_1_265;
wire    [31:0]  conv_out_1_266, conv_out_1_267, conv_out_1_268, conv_out_1_269, conv_out_1_270, conv_out_1_271, conv_out_1_272, conv_out_1_273, conv_out_1_274, conv_out_1_275, conv_out_1_276, conv_out_1_277, conv_out_1_278, conv_out_1_279;
wire    [31:0]  conv_out_1_280, conv_out_1_281, conv_out_1_282, conv_out_1_283, conv_out_1_284, conv_out_1_285, conv_out_1_286, conv_out_1_287, conv_out_1_288, conv_out_1_289, conv_out_1_290, conv_out_1_291, conv_out_1_292, conv_out_1_293;
wire    [31:0]  conv_out_1_294, conv_out_1_295, conv_out_1_296, conv_out_1_297, conv_out_1_298, conv_out_1_299, conv_out_1_300, conv_out_1_301, conv_out_1_302, conv_out_1_303, conv_out_1_304, conv_out_1_305, conv_out_1_306, conv_out_1_307;
wire    [31:0]  conv_out_1_308, conv_out_1_309, conv_out_1_310, conv_out_1_311, conv_out_1_312, conv_out_1_313, conv_out_1_314, conv_out_1_315, conv_out_1_316, conv_out_1_317, conv_out_1_318, conv_out_1_319, conv_out_1_320, conv_out_1_321;
wire    [31:0]  conv_out_1_322, conv_out_1_323, conv_out_1_324, conv_out_1_325, conv_out_1_326, conv_out_1_327, conv_out_1_328, conv_out_1_329, conv_out_1_330, conv_out_1_331, conv_out_1_332, conv_out_1_333, conv_out_1_334, conv_out_1_335;
wire    [31:0]  conv_out_1_336, conv_out_1_337, conv_out_1_338, conv_out_1_339, conv_out_1_340, conv_out_1_341, conv_out_1_342, conv_out_1_343, conv_out_1_344, conv_out_1_345, conv_out_1_346, conv_out_1_347, conv_out_1_348, conv_out_1_349;
wire    [31:0]  conv_out_1_350, conv_out_1_351, conv_out_1_352, conv_out_1_353, conv_out_1_354, conv_out_1_355, conv_out_1_356, conv_out_1_357, conv_out_1_358, conv_out_1_359, conv_out_1_360, conv_out_1_361, conv_out_1_362, conv_out_1_363;
wire    [31:0]  conv_out_1_364, conv_out_1_365, conv_out_1_366, conv_out_1_367, conv_out_1_368, conv_out_1_369, conv_out_1_370, conv_out_1_371, conv_out_1_372, conv_out_1_373, conv_out_1_374, conv_out_1_375, conv_out_1_376, conv_out_1_377;
wire    [31:0]  conv_out_1_378, conv_out_1_379, conv_out_1_380, conv_out_1_381, conv_out_1_382, conv_out_1_383, conv_out_1_384, conv_out_1_385, conv_out_1_386, conv_out_1_387, conv_out_1_388, conv_out_1_389, conv_out_1_390, conv_out_1_391;
wire    [31:0]  conv_out_1_392, conv_out_1_393, conv_out_1_394, conv_out_1_395, conv_out_1_396, conv_out_1_397, conv_out_1_398, conv_out_1_399, conv_out_1_400, conv_out_1_401, conv_out_1_402, conv_out_1_403, conv_out_1_404, conv_out_1_405;
wire    [31:0]  conv_out_1_406, conv_out_1_407, conv_out_1_408, conv_out_1_409, conv_out_1_410, conv_out_1_411, conv_out_1_412, conv_out_1_413, conv_out_1_414, conv_out_1_415, conv_out_1_416, conv_out_1_417, conv_out_1_418, conv_out_1_419;
wire    [31:0]  conv_out_1_420, conv_out_1_421, conv_out_1_422, conv_out_1_423, conv_out_1_424, conv_out_1_425, conv_out_1_426, conv_out_1_427, conv_out_1_428, conv_out_1_429, conv_out_1_430, conv_out_1_431, conv_out_1_432, conv_out_1_433;
wire    [31:0]  conv_out_1_434, conv_out_1_435, conv_out_1_436, conv_out_1_437, conv_out_1_438, conv_out_1_439, conv_out_1_440, conv_out_1_441, conv_out_1_442, conv_out_1_443, conv_out_1_444, conv_out_1_445, conv_out_1_446, conv_out_1_447;
wire    [31:0]  conv_out_1_448, conv_out_1_449, conv_out_1_450, conv_out_1_451, conv_out_1_452, conv_out_1_453, conv_out_1_454, conv_out_1_455, conv_out_1_456, conv_out_1_457, conv_out_1_458, conv_out_1_459, conv_out_1_460, conv_out_1_461;
wire    [31:0]  conv_out_1_462, conv_out_1_463, conv_out_1_464, conv_out_1_465, conv_out_1_466, conv_out_1_467, conv_out_1_468, conv_out_1_469, conv_out_1_470, conv_out_1_471, conv_out_1_472, conv_out_1_473, conv_out_1_474, conv_out_1_475;
wire    [31:0]  conv_out_1_476, conv_out_1_477, conv_out_1_478, conv_out_1_479, conv_out_1_480, conv_out_1_481, conv_out_1_482, conv_out_1_483, conv_out_1_484, conv_out_1_485, conv_out_1_486, conv_out_1_487, conv_out_1_488, conv_out_1_489;
wire    [31:0]  conv_out_1_490, conv_out_1_491, conv_out_1_492, conv_out_1_493, conv_out_1_494, conv_out_1_495, conv_out_1_496, conv_out_1_497, conv_out_1_498, conv_out_1_499, conv_out_1_500, conv_out_1_501, conv_out_1_502, conv_out_1_503;
wire    [31:0]  conv_out_1_504, conv_out_1_505, conv_out_1_506, conv_out_1_507, conv_out_1_508, conv_out_1_509, conv_out_1_510, conv_out_1_511, conv_out_1_512, conv_out_1_513, conv_out_1_514, conv_out_1_515, conv_out_1_516, conv_out_1_517;
wire    [31:0]  conv_out_1_518, conv_out_1_519, conv_out_1_520, conv_out_1_521, conv_out_1_522, conv_out_1_523, conv_out_1_524, conv_out_1_525, conv_out_1_526, conv_out_1_527, conv_out_1_528, conv_out_1_529, conv_out_1_530, conv_out_1_531;
wire    [31:0]  conv_out_1_532, conv_out_1_533, conv_out_1_534, conv_out_1_535, conv_out_1_536, conv_out_1_537, conv_out_1_538, conv_out_1_539, conv_out_1_540, conv_out_1_541, conv_out_1_542, conv_out_1_543, conv_out_1_544, conv_out_1_545;
wire    [31:0]  conv_out_1_546, conv_out_1_547, conv_out_1_548, conv_out_1_549, conv_out_1_550, conv_out_1_551, conv_out_1_552, conv_out_1_553, conv_out_1_554, conv_out_1_555, conv_out_1_556, conv_out_1_557, conv_out_1_558, conv_out_1_559;
wire    [31:0]  conv_out_1_560, conv_out_1_561, conv_out_1_562, conv_out_1_563, conv_out_1_564, conv_out_1_565, conv_out_1_566, conv_out_1_567, conv_out_1_568, conv_out_1_569, conv_out_1_570, conv_out_1_571, conv_out_1_572, conv_out_1_573;
wire    [31:0]  conv_out_1_574, conv_out_1_575, conv_out_1_576, conv_out_1_577, conv_out_1_578, conv_out_1_579, conv_out_1_580, conv_out_1_581, conv_out_1_582, conv_out_1_583, conv_out_1_584, conv_out_1_585, conv_out_1_586, conv_out_1_587;
wire    [31:0]  conv_out_1_588, conv_out_1_589, conv_out_1_590, conv_out_1_591, conv_out_1_592, conv_out_1_593, conv_out_1_594, conv_out_1_595, conv_out_1_596, conv_out_1_597, conv_out_1_598, conv_out_1_599, conv_out_1_600, conv_out_1_601;
wire    [31:0]  conv_out_1_602, conv_out_1_603, conv_out_1_604, conv_out_1_605, conv_out_1_606, conv_out_1_607, conv_out_1_608, conv_out_1_609, conv_out_1_610, conv_out_1_611, conv_out_1_612, conv_out_1_613, conv_out_1_614, conv_out_1_615;
wire    [31:0]  conv_out_1_616, conv_out_1_617, conv_out_1_618, conv_out_1_619, conv_out_1_620, conv_out_1_621, conv_out_1_622, conv_out_1_623, conv_out_1_624, conv_out_1_625, conv_out_1_626, conv_out_1_627, conv_out_1_628, conv_out_1_629;
wire    [31:0]  conv_out_1_630, conv_out_1_631, conv_out_1_632, conv_out_1_633, conv_out_1_634, conv_out_1_635, conv_out_1_636, conv_out_1_637, conv_out_1_638, conv_out_1_639, conv_out_1_640, conv_out_1_641, conv_out_1_642, conv_out_1_643;
wire    [31:0]  conv_out_1_644, conv_out_1_645, conv_out_1_646, conv_out_1_647, conv_out_1_648, conv_out_1_649, conv_out_1_650, conv_out_1_651, conv_out_1_652, conv_out_1_653, conv_out_1_654, conv_out_1_655, conv_out_1_656, conv_out_1_657;
wire    [31:0]  conv_out_1_658, conv_out_1_659, conv_out_1_660, conv_out_1_661, conv_out_1_662, conv_out_1_663, conv_out_1_664, conv_out_1_665, conv_out_1_666, conv_out_1_667, conv_out_1_668, conv_out_1_669, conv_out_1_670, conv_out_1_671;
wire    [31:0]  conv_out_1_672, conv_out_1_673, conv_out_1_674, conv_out_1_675, conv_out_1_676, conv_out_1_677, conv_out_1_678, conv_out_1_679, conv_out_1_680, conv_out_1_681, conv_out_1_682, conv_out_1_683, conv_out_1_684, conv_out_1_685;
wire    [31:0]  conv_out_1_686, conv_out_1_687, conv_out_1_688, conv_out_1_689, conv_out_1_690, conv_out_1_691, conv_out_1_692, conv_out_1_693, conv_out_1_694, conv_out_1_695, conv_out_1_696, conv_out_1_697, conv_out_1_698, conv_out_1_699;
wire    [31:0]  conv_out_1_700, conv_out_1_701, conv_out_1_702, conv_out_1_703, conv_out_1_704, conv_out_1_705, conv_out_1_706, conv_out_1_707, conv_out_1_708, conv_out_1_709, conv_out_1_710, conv_out_1_711, conv_out_1_712, conv_out_1_713;
wire    [31:0]  conv_out_1_714, conv_out_1_715, conv_out_1_716, conv_out_1_717, conv_out_1_718, conv_out_1_719, conv_out_1_720, conv_out_1_721, conv_out_1_722, conv_out_1_723, conv_out_1_724, conv_out_1_725, conv_out_1_726, conv_out_1_727;
wire    [31:0]  conv_out_1_728, conv_out_1_729, conv_out_1_730, conv_out_1_731, conv_out_1_732, conv_out_1_733, conv_out_1_734, conv_out_1_735, conv_out_1_736, conv_out_1_737, conv_out_1_738, conv_out_1_739, conv_out_1_740, conv_out_1_741;
wire    [31:0]  conv_out_1_742, conv_out_1_743, conv_out_1_744, conv_out_1_745, conv_out_1_746, conv_out_1_747, conv_out_1_748, conv_out_1_749, conv_out_1_750, conv_out_1_751, conv_out_1_752, conv_out_1_753, conv_out_1_754, conv_out_1_755;
wire    [31:0]  conv_out_1_756, conv_out_1_757, conv_out_1_758, conv_out_1_759, conv_out_1_760, conv_out_1_761, conv_out_1_762, conv_out_1_763, conv_out_1_764, conv_out_1_765, conv_out_1_766, conv_out_1_767, conv_out_1_768, conv_out_1_769;
wire    [31:0]  conv_out_1_770, conv_out_1_771, conv_out_1_772, conv_out_1_773, conv_out_1_774, conv_out_1_775, conv_out_1_776, conv_out_1_777, conv_out_1_778, conv_out_1_779, conv_out_1_780, conv_out_1_781, conv_out_1_782, conv_out_1_783;

    assign  image_1_0[143:128]   = Conv_out[899];
    assign  image_1_0[127:112]   = Conv_out[898];
    assign  image_1_0[111:96]    = Conv_out[897];
    assign  image_1_0[95:80]     = Conv_out[869];
    assign  image_1_0[79:64]     = Conv_out[868];
    assign  image_1_0[63:48]     = Conv_out[867];
    assign  image_1_0[47:32]     = Conv_out[839];
    assign  image_1_0[31:16]     = Conv_out[838];
    assign  image_1_0[15:0]      = Conv_out[837];

    assign  image_1_1[143:128]   = Conv_out[898];
    assign  image_1_1[127:112]   = Conv_out[897];
    assign  image_1_1[111:96]    = Conv_out[896];
    assign  image_1_1[95:80]     = Conv_out[868];
    assign  image_1_1[79:64]     = Conv_out[867];
    assign  image_1_1[63:48]     = Conv_out[866];
    assign  image_1_1[47:32]     = Conv_out[838];
    assign  image_1_1[31:16]     = Conv_out[837];
    assign  image_1_1[15:0]      = Conv_out[836];

    assign  image_1_2[143:128]   = Conv_out[897];
    assign  image_1_2[127:112]   = Conv_out[896];
    assign  image_1_2[111:96]    = Conv_out[895];
    assign  image_1_2[95:80]     = Conv_out[867];
    assign  image_1_2[79:64]     = Conv_out[866];
    assign  image_1_2[63:48]     = Conv_out[865];
    assign  image_1_2[47:32]     = Conv_out[837];
    assign  image_1_2[31:16]     = Conv_out[836];
    assign  image_1_2[15:0]      = Conv_out[835];

    assign  image_1_3[143:128]   = Conv_out[896];
    assign  image_1_3[127:112]   = Conv_out[895];
    assign  image_1_3[111:96]    = Conv_out[894];
    assign  image_1_3[95:80]     = Conv_out[866];
    assign  image_1_3[79:64]     = Conv_out[865];
    assign  image_1_3[63:48]     = Conv_out[864];
    assign  image_1_3[47:32]     = Conv_out[836];
    assign  image_1_3[31:16]     = Conv_out[835];
    assign  image_1_3[15:0]      = Conv_out[834];

    assign  image_1_4[143:128]   = Conv_out[895];
    assign  image_1_4[127:112]   = Conv_out[894];
    assign  image_1_4[111:96]    = Conv_out[893];
    assign  image_1_4[95:80]     = Conv_out[865];
    assign  image_1_4[79:64]     = Conv_out[864];
    assign  image_1_4[63:48]     = Conv_out[863];
    assign  image_1_4[47:32]     = Conv_out[835];
    assign  image_1_4[31:16]     = Conv_out[834];
    assign  image_1_4[15:0]      = Conv_out[833];

    assign  image_1_5[143:128]   = Conv_out[894];
    assign  image_1_5[127:112]   = Conv_out[893];
    assign  image_1_5[111:96]    = Conv_out[892];
    assign  image_1_5[95:80]     = Conv_out[864];
    assign  image_1_5[79:64]     = Conv_out[863];
    assign  image_1_5[63:48]     = Conv_out[862];
    assign  image_1_5[47:32]     = Conv_out[834];
    assign  image_1_5[31:16]     = Conv_out[833];
    assign  image_1_5[15:0]      = Conv_out[832];

    assign  image_1_6[143:128]   = Conv_out[893];
    assign  image_1_6[127:112]   = Conv_out[892];
    assign  image_1_6[111:96]    = Conv_out[891];
    assign  image_1_6[95:80]     = Conv_out[863];
    assign  image_1_6[79:64]     = Conv_out[862];
    assign  image_1_6[63:48]     = Conv_out[861];
    assign  image_1_6[47:32]     = Conv_out[833];
    assign  image_1_6[31:16]     = Conv_out[832];
    assign  image_1_6[15:0]      = Conv_out[831];

    assign  image_1_7[143:128]   = Conv_out[892];
    assign  image_1_7[127:112]   = Conv_out[891];
    assign  image_1_7[111:96]    = Conv_out[890];
    assign  image_1_7[95:80]     = Conv_out[862];
    assign  image_1_7[79:64]     = Conv_out[861];
    assign  image_1_7[63:48]     = Conv_out[860];
    assign  image_1_7[47:32]     = Conv_out[832];
    assign  image_1_7[31:16]     = Conv_out[831];
    assign  image_1_7[15:0]      = Conv_out[830];

    assign  image_1_8[143:128]   = Conv_out[891];
    assign  image_1_8[127:112]   = Conv_out[890];
    assign  image_1_8[111:96]    = Conv_out[889];
    assign  image_1_8[95:80]     = Conv_out[861];
    assign  image_1_8[79:64]     = Conv_out[860];
    assign  image_1_8[63:48]     = Conv_out[859];
    assign  image_1_8[47:32]     = Conv_out[831];
    assign  image_1_8[31:16]     = Conv_out[830];
    assign  image_1_8[15:0]      = Conv_out[829];

    assign  image_1_9[143:128]   = Conv_out[890];
    assign  image_1_9[127:112]   = Conv_out[889];
    assign  image_1_9[111:96]    = Conv_out[888];
    assign  image_1_9[95:80]     = Conv_out[860];
    assign  image_1_9[79:64]     = Conv_out[859];
    assign  image_1_9[63:48]     = Conv_out[858];
    assign  image_1_9[47:32]     = Conv_out[830];
    assign  image_1_9[31:16]     = Conv_out[829];
    assign  image_1_9[15:0]      = Conv_out[828];

    assign  image_1_10[143:128]   = Conv_out[889];
    assign  image_1_10[127:112]   = Conv_out[888];
    assign  image_1_10[111:96]    = Conv_out[887];
    assign  image_1_10[95:80]     = Conv_out[859];
    assign  image_1_10[79:64]     = Conv_out[858];
    assign  image_1_10[63:48]     = Conv_out[857];
    assign  image_1_10[47:32]     = Conv_out[829];
    assign  image_1_10[31:16]     = Conv_out[828];
    assign  image_1_10[15:0]      = Conv_out[827];

    assign  image_1_11[143:128]   = Conv_out[888];
    assign  image_1_11[127:112]   = Conv_out[887];
    assign  image_1_11[111:96]    = Conv_out[886];
    assign  image_1_11[95:80]     = Conv_out[858];
    assign  image_1_11[79:64]     = Conv_out[857];
    assign  image_1_11[63:48]     = Conv_out[856];
    assign  image_1_11[47:32]     = Conv_out[828];
    assign  image_1_11[31:16]     = Conv_out[827];
    assign  image_1_11[15:0]      = Conv_out[826];

    assign  image_1_12[143:128]   = Conv_out[887];
    assign  image_1_12[127:112]   = Conv_out[886];
    assign  image_1_12[111:96]    = Conv_out[885];
    assign  image_1_12[95:80]     = Conv_out[857];
    assign  image_1_12[79:64]     = Conv_out[856];
    assign  image_1_12[63:48]     = Conv_out[855];
    assign  image_1_12[47:32]     = Conv_out[827];
    assign  image_1_12[31:16]     = Conv_out[826];
    assign  image_1_12[15:0]      = Conv_out[825];

    assign  image_1_13[143:128]   = Conv_out[886];
    assign  image_1_13[127:112]   = Conv_out[885];
    assign  image_1_13[111:96]    = Conv_out[884];
    assign  image_1_13[95:80]     = Conv_out[856];
    assign  image_1_13[79:64]     = Conv_out[855];
    assign  image_1_13[63:48]     = Conv_out[854];
    assign  image_1_13[47:32]     = Conv_out[826];
    assign  image_1_13[31:16]     = Conv_out[825];
    assign  image_1_13[15:0]      = Conv_out[824];

    assign  image_1_14[143:128]   = Conv_out[885];
    assign  image_1_14[127:112]   = Conv_out[884];
    assign  image_1_14[111:96]    = Conv_out[883];
    assign  image_1_14[95:80]     = Conv_out[855];
    assign  image_1_14[79:64]     = Conv_out[854];
    assign  image_1_14[63:48]     = Conv_out[853];
    assign  image_1_14[47:32]     = Conv_out[825];
    assign  image_1_14[31:16]     = Conv_out[824];
    assign  image_1_14[15:0]      = Conv_out[823];

    assign  image_1_15[143:128]   = Conv_out[884];
    assign  image_1_15[127:112]   = Conv_out[883];
    assign  image_1_15[111:96]    = Conv_out[882];
    assign  image_1_15[95:80]     = Conv_out[854];
    assign  image_1_15[79:64]     = Conv_out[853];
    assign  image_1_15[63:48]     = Conv_out[852];
    assign  image_1_15[47:32]     = Conv_out[824];
    assign  image_1_15[31:16]     = Conv_out[823];
    assign  image_1_15[15:0]      = Conv_out[822];

    assign  image_1_16[143:128]   = Conv_out[883];
    assign  image_1_16[127:112]   = Conv_out[882];
    assign  image_1_16[111:96]    = Conv_out[881];
    assign  image_1_16[95:80]     = Conv_out[853];
    assign  image_1_16[79:64]     = Conv_out[852];
    assign  image_1_16[63:48]     = Conv_out[851];
    assign  image_1_16[47:32]     = Conv_out[823];
    assign  image_1_16[31:16]     = Conv_out[822];
    assign  image_1_16[15:0]      = Conv_out[821];

    assign  image_1_17[143:128]   = Conv_out[882];
    assign  image_1_17[127:112]   = Conv_out[881];
    assign  image_1_17[111:96]    = Conv_out[880];
    assign  image_1_17[95:80]     = Conv_out[852];
    assign  image_1_17[79:64]     = Conv_out[851];
    assign  image_1_17[63:48]     = Conv_out[850];
    assign  image_1_17[47:32]     = Conv_out[822];
    assign  image_1_17[31:16]     = Conv_out[821];
    assign  image_1_17[15:0]      = Conv_out[820];

    assign  image_1_18[143:128]   = Conv_out[881];
    assign  image_1_18[127:112]   = Conv_out[880];
    assign  image_1_18[111:96]    = Conv_out[879];
    assign  image_1_18[95:80]     = Conv_out[851];
    assign  image_1_18[79:64]     = Conv_out[850];
    assign  image_1_18[63:48]     = Conv_out[849];
    assign  image_1_18[47:32]     = Conv_out[821];
    assign  image_1_18[31:16]     = Conv_out[820];
    assign  image_1_18[15:0]      = Conv_out[819];

    assign  image_1_19[143:128]   = Conv_out[880];
    assign  image_1_19[127:112]   = Conv_out[879];
    assign  image_1_19[111:96]    = Conv_out[878];
    assign  image_1_19[95:80]     = Conv_out[850];
    assign  image_1_19[79:64]     = Conv_out[849];
    assign  image_1_19[63:48]     = Conv_out[848];
    assign  image_1_19[47:32]     = Conv_out[820];
    assign  image_1_19[31:16]     = Conv_out[819];
    assign  image_1_19[15:0]      = Conv_out[818];

    assign  image_1_20[143:128]   = Conv_out[879];
    assign  image_1_20[127:112]   = Conv_out[878];
    assign  image_1_20[111:96]    = Conv_out[877];
    assign  image_1_20[95:80]     = Conv_out[849];
    assign  image_1_20[79:64]     = Conv_out[848];
    assign  image_1_20[63:48]     = Conv_out[847];
    assign  image_1_20[47:32]     = Conv_out[819];
    assign  image_1_20[31:16]     = Conv_out[818];
    assign  image_1_20[15:0]      = Conv_out[817];

    assign  image_1_21[143:128]   = Conv_out[878];
    assign  image_1_21[127:112]   = Conv_out[877];
    assign  image_1_21[111:96]    = Conv_out[876];
    assign  image_1_21[95:80]     = Conv_out[848];
    assign  image_1_21[79:64]     = Conv_out[847];
    assign  image_1_21[63:48]     = Conv_out[846];
    assign  image_1_21[47:32]     = Conv_out[818];
    assign  image_1_21[31:16]     = Conv_out[817];
    assign  image_1_21[15:0]      = Conv_out[816];

    assign  image_1_22[143:128]   = Conv_out[877];
    assign  image_1_22[127:112]   = Conv_out[876];
    assign  image_1_22[111:96]    = Conv_out[875];
    assign  image_1_22[95:80]     = Conv_out[847];
    assign  image_1_22[79:64]     = Conv_out[846];
    assign  image_1_22[63:48]     = Conv_out[845];
    assign  image_1_22[47:32]     = Conv_out[817];
    assign  image_1_22[31:16]     = Conv_out[816];
    assign  image_1_22[15:0]      = Conv_out[815];

    assign  image_1_23[143:128]   = Conv_out[876];
    assign  image_1_23[127:112]   = Conv_out[875];
    assign  image_1_23[111:96]    = Conv_out[874];
    assign  image_1_23[95:80]     = Conv_out[846];
    assign  image_1_23[79:64]     = Conv_out[845];
    assign  image_1_23[63:48]     = Conv_out[844];
    assign  image_1_23[47:32]     = Conv_out[816];
    assign  image_1_23[31:16]     = Conv_out[815];
    assign  image_1_23[15:0]      = Conv_out[814];

    assign  image_1_24[143:128]   = Conv_out[875];
    assign  image_1_24[127:112]   = Conv_out[874];
    assign  image_1_24[111:96]    = Conv_out[873];
    assign  image_1_24[95:80]     = Conv_out[845];
    assign  image_1_24[79:64]     = Conv_out[844];
    assign  image_1_24[63:48]     = Conv_out[843];
    assign  image_1_24[47:32]     = Conv_out[815];
    assign  image_1_24[31:16]     = Conv_out[814];
    assign  image_1_24[15:0]      = Conv_out[813];

    assign  image_1_25[143:128]   = Conv_out[874];
    assign  image_1_25[127:112]   = Conv_out[873];
    assign  image_1_25[111:96]    = Conv_out[872];
    assign  image_1_25[95:80]     = Conv_out[844];
    assign  image_1_25[79:64]     = Conv_out[843];
    assign  image_1_25[63:48]     = Conv_out[842];
    assign  image_1_25[47:32]     = Conv_out[814];
    assign  image_1_25[31:16]     = Conv_out[813];
    assign  image_1_25[15:0]      = Conv_out[812];

    assign  image_1_26[143:128]   = Conv_out[873];
    assign  image_1_26[127:112]   = Conv_out[872];
    assign  image_1_26[111:96]    = Conv_out[871];
    assign  image_1_26[95:80]     = Conv_out[843];
    assign  image_1_26[79:64]     = Conv_out[842];
    assign  image_1_26[63:48]     = Conv_out[841];
    assign  image_1_26[47:32]     = Conv_out[813];
    assign  image_1_26[31:16]     = Conv_out[812];
    assign  image_1_26[15:0]      = Conv_out[811];

    assign  image_1_27[143:128]   = Conv_out[872];
    assign  image_1_27[127:112]   = Conv_out[871];
    assign  image_1_27[111:96]    = Conv_out[870];
    assign  image_1_27[95:80]     = Conv_out[842];
    assign  image_1_27[79:64]     = Conv_out[841];
    assign  image_1_27[63:48]     = Conv_out[840];
    assign  image_1_27[47:32]     = Conv_out[812];
    assign  image_1_27[31:16]     = Conv_out[811];
    assign  image_1_27[15:0]      = Conv_out[810];

    assign  image_1_28[143:128]   = Conv_out[869];
    assign  image_1_28[127:112]   = Conv_out[868];
    assign  image_1_28[111:96]    = Conv_out[867];
    assign  image_1_28[95:80]     = Conv_out[839];
    assign  image_1_28[79:64]     = Conv_out[838];
    assign  image_1_28[63:48]     = Conv_out[837];
    assign  image_1_28[47:32]     = Conv_out[809];
    assign  image_1_28[31:16]     = Conv_out[808];
    assign  image_1_28[15:0]      = Conv_out[807];

    assign  image_1_29[143:128]   = Conv_out[868];
    assign  image_1_29[127:112]   = Conv_out[867];
    assign  image_1_29[111:96]    = Conv_out[866];
    assign  image_1_29[95:80]     = Conv_out[838];
    assign  image_1_29[79:64]     = Conv_out[837];
    assign  image_1_29[63:48]     = Conv_out[836];
    assign  image_1_29[47:32]     = Conv_out[808];
    assign  image_1_29[31:16]     = Conv_out[807];
    assign  image_1_29[15:0]      = Conv_out[806];

    assign  image_1_30[143:128]   = Conv_out[867];
    assign  image_1_30[127:112]   = Conv_out[866];
    assign  image_1_30[111:96]    = Conv_out[865];
    assign  image_1_30[95:80]     = Conv_out[837];
    assign  image_1_30[79:64]     = Conv_out[836];
    assign  image_1_30[63:48]     = Conv_out[835];
    assign  image_1_30[47:32]     = Conv_out[807];
    assign  image_1_30[31:16]     = Conv_out[806];
    assign  image_1_30[15:0]      = Conv_out[805];

    assign  image_1_31[143:128]   = Conv_out[866];
    assign  image_1_31[127:112]   = Conv_out[865];
    assign  image_1_31[111:96]    = Conv_out[864];
    assign  image_1_31[95:80]     = Conv_out[836];
    assign  image_1_31[79:64]     = Conv_out[835];
    assign  image_1_31[63:48]     = Conv_out[834];
    assign  image_1_31[47:32]     = Conv_out[806];
    assign  image_1_31[31:16]     = Conv_out[805];
    assign  image_1_31[15:0]      = Conv_out[804];

    assign  image_1_32[143:128]   = Conv_out[865];
    assign  image_1_32[127:112]   = Conv_out[864];
    assign  image_1_32[111:96]    = Conv_out[863];
    assign  image_1_32[95:80]     = Conv_out[835];
    assign  image_1_32[79:64]     = Conv_out[834];
    assign  image_1_32[63:48]     = Conv_out[833];
    assign  image_1_32[47:32]     = Conv_out[805];
    assign  image_1_32[31:16]     = Conv_out[804];
    assign  image_1_32[15:0]      = Conv_out[803];

    assign  image_1_33[143:128]   = Conv_out[864];
    assign  image_1_33[127:112]   = Conv_out[863];
    assign  image_1_33[111:96]    = Conv_out[862];
    assign  image_1_33[95:80]     = Conv_out[834];
    assign  image_1_33[79:64]     = Conv_out[833];
    assign  image_1_33[63:48]     = Conv_out[832];
    assign  image_1_33[47:32]     = Conv_out[804];
    assign  image_1_33[31:16]     = Conv_out[803];
    assign  image_1_33[15:0]      = Conv_out[802];

    assign  image_1_34[143:128]   = Conv_out[863];
    assign  image_1_34[127:112]   = Conv_out[862];
    assign  image_1_34[111:96]    = Conv_out[861];
    assign  image_1_34[95:80]     = Conv_out[833];
    assign  image_1_34[79:64]     = Conv_out[832];
    assign  image_1_34[63:48]     = Conv_out[831];
    assign  image_1_34[47:32]     = Conv_out[803];
    assign  image_1_34[31:16]     = Conv_out[802];
    assign  image_1_34[15:0]      = Conv_out[801];

    assign  image_1_35[143:128]   = Conv_out[862];
    assign  image_1_35[127:112]   = Conv_out[861];
    assign  image_1_35[111:96]    = Conv_out[860];
    assign  image_1_35[95:80]     = Conv_out[832];
    assign  image_1_35[79:64]     = Conv_out[831];
    assign  image_1_35[63:48]     = Conv_out[830];
    assign  image_1_35[47:32]     = Conv_out[802];
    assign  image_1_35[31:16]     = Conv_out[801];
    assign  image_1_35[15:0]      = Conv_out[800];

    assign  image_1_36[143:128]   = Conv_out[861];
    assign  image_1_36[127:112]   = Conv_out[860];
    assign  image_1_36[111:96]    = Conv_out[859];
    assign  image_1_36[95:80]     = Conv_out[831];
    assign  image_1_36[79:64]     = Conv_out[830];
    assign  image_1_36[63:48]     = Conv_out[829];
    assign  image_1_36[47:32]     = Conv_out[801];
    assign  image_1_36[31:16]     = Conv_out[800];
    assign  image_1_36[15:0]      = Conv_out[799];

    assign  image_1_37[143:128]   = Conv_out[860];
    assign  image_1_37[127:112]   = Conv_out[859];
    assign  image_1_37[111:96]    = Conv_out[858];
    assign  image_1_37[95:80]     = Conv_out[830];
    assign  image_1_37[79:64]     = Conv_out[829];
    assign  image_1_37[63:48]     = Conv_out[828];
    assign  image_1_37[47:32]     = Conv_out[800];
    assign  image_1_37[31:16]     = Conv_out[799];
    assign  image_1_37[15:0]      = Conv_out[798];

    assign  image_1_38[143:128]   = Conv_out[859];
    assign  image_1_38[127:112]   = Conv_out[858];
    assign  image_1_38[111:96]    = Conv_out[857];
    assign  image_1_38[95:80]     = Conv_out[829];
    assign  image_1_38[79:64]     = Conv_out[828];
    assign  image_1_38[63:48]     = Conv_out[827];
    assign  image_1_38[47:32]     = Conv_out[799];
    assign  image_1_38[31:16]     = Conv_out[798];
    assign  image_1_38[15:0]      = Conv_out[797];

    assign  image_1_39[143:128]   = Conv_out[858];
    assign  image_1_39[127:112]   = Conv_out[857];
    assign  image_1_39[111:96]    = Conv_out[856];
    assign  image_1_39[95:80]     = Conv_out[828];
    assign  image_1_39[79:64]     = Conv_out[827];
    assign  image_1_39[63:48]     = Conv_out[826];
    assign  image_1_39[47:32]     = Conv_out[798];
    assign  image_1_39[31:16]     = Conv_out[797];
    assign  image_1_39[15:0]      = Conv_out[796];

    assign  image_1_40[143:128]   = Conv_out[857];
    assign  image_1_40[127:112]   = Conv_out[856];
    assign  image_1_40[111:96]    = Conv_out[855];
    assign  image_1_40[95:80]     = Conv_out[827];
    assign  image_1_40[79:64]     = Conv_out[826];
    assign  image_1_40[63:48]     = Conv_out[825];
    assign  image_1_40[47:32]     = Conv_out[797];
    assign  image_1_40[31:16]     = Conv_out[796];
    assign  image_1_40[15:0]      = Conv_out[795];

    assign  image_1_41[143:128]   = Conv_out[856];
    assign  image_1_41[127:112]   = Conv_out[855];
    assign  image_1_41[111:96]    = Conv_out[854];
    assign  image_1_41[95:80]     = Conv_out[826];
    assign  image_1_41[79:64]     = Conv_out[825];
    assign  image_1_41[63:48]     = Conv_out[824];
    assign  image_1_41[47:32]     = Conv_out[796];
    assign  image_1_41[31:16]     = Conv_out[795];
    assign  image_1_41[15:0]      = Conv_out[794];

    assign  image_1_42[143:128]   = Conv_out[855];
    assign  image_1_42[127:112]   = Conv_out[854];
    assign  image_1_42[111:96]    = Conv_out[853];
    assign  image_1_42[95:80]     = Conv_out[825];
    assign  image_1_42[79:64]     = Conv_out[824];
    assign  image_1_42[63:48]     = Conv_out[823];
    assign  image_1_42[47:32]     = Conv_out[795];
    assign  image_1_42[31:16]     = Conv_out[794];
    assign  image_1_42[15:0]      = Conv_out[793];

    assign  image_1_43[143:128]   = Conv_out[854];
    assign  image_1_43[127:112]   = Conv_out[853];
    assign  image_1_43[111:96]    = Conv_out[852];
    assign  image_1_43[95:80]     = Conv_out[824];
    assign  image_1_43[79:64]     = Conv_out[823];
    assign  image_1_43[63:48]     = Conv_out[822];
    assign  image_1_43[47:32]     = Conv_out[794];
    assign  image_1_43[31:16]     = Conv_out[793];
    assign  image_1_43[15:0]      = Conv_out[792];

    assign  image_1_44[143:128]   = Conv_out[853];
    assign  image_1_44[127:112]   = Conv_out[852];
    assign  image_1_44[111:96]    = Conv_out[851];
    assign  image_1_44[95:80]     = Conv_out[823];
    assign  image_1_44[79:64]     = Conv_out[822];
    assign  image_1_44[63:48]     = Conv_out[821];
    assign  image_1_44[47:32]     = Conv_out[793];
    assign  image_1_44[31:16]     = Conv_out[792];
    assign  image_1_44[15:0]      = Conv_out[791];

    assign  image_1_45[143:128]   = Conv_out[852];
    assign  image_1_45[127:112]   = Conv_out[851];
    assign  image_1_45[111:96]    = Conv_out[850];
    assign  image_1_45[95:80]     = Conv_out[822];
    assign  image_1_45[79:64]     = Conv_out[821];
    assign  image_1_45[63:48]     = Conv_out[820];
    assign  image_1_45[47:32]     = Conv_out[792];
    assign  image_1_45[31:16]     = Conv_out[791];
    assign  image_1_45[15:0]      = Conv_out[790];

    assign  image_1_46[143:128]   = Conv_out[851];
    assign  image_1_46[127:112]   = Conv_out[850];
    assign  image_1_46[111:96]    = Conv_out[849];
    assign  image_1_46[95:80]     = Conv_out[821];
    assign  image_1_46[79:64]     = Conv_out[820];
    assign  image_1_46[63:48]     = Conv_out[819];
    assign  image_1_46[47:32]     = Conv_out[791];
    assign  image_1_46[31:16]     = Conv_out[790];
    assign  image_1_46[15:0]      = Conv_out[789];

    assign  image_1_47[143:128]   = Conv_out[850];
    assign  image_1_47[127:112]   = Conv_out[849];
    assign  image_1_47[111:96]    = Conv_out[848];
    assign  image_1_47[95:80]     = Conv_out[820];
    assign  image_1_47[79:64]     = Conv_out[819];
    assign  image_1_47[63:48]     = Conv_out[818];
    assign  image_1_47[47:32]     = Conv_out[790];
    assign  image_1_47[31:16]     = Conv_out[789];
    assign  image_1_47[15:0]      = Conv_out[788];

    assign  image_1_48[143:128]   = Conv_out[849];
    assign  image_1_48[127:112]   = Conv_out[848];
    assign  image_1_48[111:96]    = Conv_out[847];
    assign  image_1_48[95:80]     = Conv_out[819];
    assign  image_1_48[79:64]     = Conv_out[818];
    assign  image_1_48[63:48]     = Conv_out[817];
    assign  image_1_48[47:32]     = Conv_out[789];
    assign  image_1_48[31:16]     = Conv_out[788];
    assign  image_1_48[15:0]      = Conv_out[787];

    assign  image_1_49[143:128]   = Conv_out[848];
    assign  image_1_49[127:112]   = Conv_out[847];
    assign  image_1_49[111:96]    = Conv_out[846];
    assign  image_1_49[95:80]     = Conv_out[818];
    assign  image_1_49[79:64]     = Conv_out[817];
    assign  image_1_49[63:48]     = Conv_out[816];
    assign  image_1_49[47:32]     = Conv_out[788];
    assign  image_1_49[31:16]     = Conv_out[787];
    assign  image_1_49[15:0]      = Conv_out[786];

    assign  image_1_50[143:128]   = Conv_out[847];
    assign  image_1_50[127:112]   = Conv_out[846];
    assign  image_1_50[111:96]    = Conv_out[845];
    assign  image_1_50[95:80]     = Conv_out[817];
    assign  image_1_50[79:64]     = Conv_out[816];
    assign  image_1_50[63:48]     = Conv_out[815];
    assign  image_1_50[47:32]     = Conv_out[787];
    assign  image_1_50[31:16]     = Conv_out[786];
    assign  image_1_50[15:0]      = Conv_out[785];

    assign  image_1_51[143:128]   = Conv_out[846];
    assign  image_1_51[127:112]   = Conv_out[845];
    assign  image_1_51[111:96]    = Conv_out[844];
    assign  image_1_51[95:80]     = Conv_out[816];
    assign  image_1_51[79:64]     = Conv_out[815];
    assign  image_1_51[63:48]     = Conv_out[814];
    assign  image_1_51[47:32]     = Conv_out[786];
    assign  image_1_51[31:16]     = Conv_out[785];
    assign  image_1_51[15:0]      = Conv_out[784];

    assign  image_1_52[143:128]   = Conv_out[845];
    assign  image_1_52[127:112]   = Conv_out[844];
    assign  image_1_52[111:96]    = Conv_out[843];
    assign  image_1_52[95:80]     = Conv_out[815];
    assign  image_1_52[79:64]     = Conv_out[814];
    assign  image_1_52[63:48]     = Conv_out[813];
    assign  image_1_52[47:32]     = Conv_out[785];
    assign  image_1_52[31:16]     = Conv_out[784];
    assign  image_1_52[15:0]      = Conv_out[783];

    assign  image_1_53[143:128]   = Conv_out[844];
    assign  image_1_53[127:112]   = Conv_out[843];
    assign  image_1_53[111:96]    = Conv_out[842];
    assign  image_1_53[95:80]     = Conv_out[814];
    assign  image_1_53[79:64]     = Conv_out[813];
    assign  image_1_53[63:48]     = Conv_out[812];
    assign  image_1_53[47:32]     = Conv_out[784];
    assign  image_1_53[31:16]     = Conv_out[783];
    assign  image_1_53[15:0]      = Conv_out[782];

    assign  image_1_54[143:128]   = Conv_out[843];
    assign  image_1_54[127:112]   = Conv_out[842];
    assign  image_1_54[111:96]    = Conv_out[841];
    assign  image_1_54[95:80]     = Conv_out[813];
    assign  image_1_54[79:64]     = Conv_out[812];
    assign  image_1_54[63:48]     = Conv_out[811];
    assign  image_1_54[47:32]     = Conv_out[783];
    assign  image_1_54[31:16]     = Conv_out[782];
    assign  image_1_54[15:0]      = Conv_out[781];

    assign  image_1_55[143:128]   = Conv_out[842];
    assign  image_1_55[127:112]   = Conv_out[841];
    assign  image_1_55[111:96]    = Conv_out[840];
    assign  image_1_55[95:80]     = Conv_out[812];
    assign  image_1_55[79:64]     = Conv_out[811];
    assign  image_1_55[63:48]     = Conv_out[810];
    assign  image_1_55[47:32]     = Conv_out[782];
    assign  image_1_55[31:16]     = Conv_out[781];
    assign  image_1_55[15:0]      = Conv_out[780];

    assign  image_1_56[143:128]   = Conv_out[839];
    assign  image_1_56[127:112]   = Conv_out[838];
    assign  image_1_56[111:96]    = Conv_out[837];
    assign  image_1_56[95:80]     = Conv_out[809];
    assign  image_1_56[79:64]     = Conv_out[808];
    assign  image_1_56[63:48]     = Conv_out[807];
    assign  image_1_56[47:32]     = Conv_out[779];
    assign  image_1_56[31:16]     = Conv_out[778];
    assign  image_1_56[15:0]      = Conv_out[777];

    assign  image_1_57[143:128]   = Conv_out[838];
    assign  image_1_57[127:112]   = Conv_out[837];
    assign  image_1_57[111:96]    = Conv_out[836];
    assign  image_1_57[95:80]     = Conv_out[808];
    assign  image_1_57[79:64]     = Conv_out[807];
    assign  image_1_57[63:48]     = Conv_out[806];
    assign  image_1_57[47:32]     = Conv_out[778];
    assign  image_1_57[31:16]     = Conv_out[777];
    assign  image_1_57[15:0]      = Conv_out[776];

    assign  image_1_58[143:128]   = Conv_out[837];
    assign  image_1_58[127:112]   = Conv_out[836];
    assign  image_1_58[111:96]    = Conv_out[835];
    assign  image_1_58[95:80]     = Conv_out[807];
    assign  image_1_58[79:64]     = Conv_out[806];
    assign  image_1_58[63:48]     = Conv_out[805];
    assign  image_1_58[47:32]     = Conv_out[777];
    assign  image_1_58[31:16]     = Conv_out[776];
    assign  image_1_58[15:0]      = Conv_out[775];

    assign  image_1_59[143:128]   = Conv_out[836];
    assign  image_1_59[127:112]   = Conv_out[835];
    assign  image_1_59[111:96]    = Conv_out[834];
    assign  image_1_59[95:80]     = Conv_out[806];
    assign  image_1_59[79:64]     = Conv_out[805];
    assign  image_1_59[63:48]     = Conv_out[804];
    assign  image_1_59[47:32]     = Conv_out[776];
    assign  image_1_59[31:16]     = Conv_out[775];
    assign  image_1_59[15:0]      = Conv_out[774];

    assign  image_1_60[143:128]   = Conv_out[835];
    assign  image_1_60[127:112]   = Conv_out[834];
    assign  image_1_60[111:96]    = Conv_out[833];
    assign  image_1_60[95:80]     = Conv_out[805];
    assign  image_1_60[79:64]     = Conv_out[804];
    assign  image_1_60[63:48]     = Conv_out[803];
    assign  image_1_60[47:32]     = Conv_out[775];
    assign  image_1_60[31:16]     = Conv_out[774];
    assign  image_1_60[15:0]      = Conv_out[773];

    assign  image_1_61[143:128]   = Conv_out[834];
    assign  image_1_61[127:112]   = Conv_out[833];
    assign  image_1_61[111:96]    = Conv_out[832];
    assign  image_1_61[95:80]     = Conv_out[804];
    assign  image_1_61[79:64]     = Conv_out[803];
    assign  image_1_61[63:48]     = Conv_out[802];
    assign  image_1_61[47:32]     = Conv_out[774];
    assign  image_1_61[31:16]     = Conv_out[773];
    assign  image_1_61[15:0]      = Conv_out[772];

    assign  image_1_62[143:128]   = Conv_out[833];
    assign  image_1_62[127:112]   = Conv_out[832];
    assign  image_1_62[111:96]    = Conv_out[831];
    assign  image_1_62[95:80]     = Conv_out[803];
    assign  image_1_62[79:64]     = Conv_out[802];
    assign  image_1_62[63:48]     = Conv_out[801];
    assign  image_1_62[47:32]     = Conv_out[773];
    assign  image_1_62[31:16]     = Conv_out[772];
    assign  image_1_62[15:0]      = Conv_out[771];

    assign  image_1_63[143:128]   = Conv_out[832];
    assign  image_1_63[127:112]   = Conv_out[831];
    assign  image_1_63[111:96]    = Conv_out[830];
    assign  image_1_63[95:80]     = Conv_out[802];
    assign  image_1_63[79:64]     = Conv_out[801];
    assign  image_1_63[63:48]     = Conv_out[800];
    assign  image_1_63[47:32]     = Conv_out[772];
    assign  image_1_63[31:16]     = Conv_out[771];
    assign  image_1_63[15:0]      = Conv_out[770];

    assign  image_1_64[143:128]   = Conv_out[831];
    assign  image_1_64[127:112]   = Conv_out[830];
    assign  image_1_64[111:96]    = Conv_out[829];
    assign  image_1_64[95:80]     = Conv_out[801];
    assign  image_1_64[79:64]     = Conv_out[800];
    assign  image_1_64[63:48]     = Conv_out[799];
    assign  image_1_64[47:32]     = Conv_out[771];
    assign  image_1_64[31:16]     = Conv_out[770];
    assign  image_1_64[15:0]      = Conv_out[769];

    assign  image_1_65[143:128]   = Conv_out[830];
    assign  image_1_65[127:112]   = Conv_out[829];
    assign  image_1_65[111:96]    = Conv_out[828];
    assign  image_1_65[95:80]     = Conv_out[800];
    assign  image_1_65[79:64]     = Conv_out[799];
    assign  image_1_65[63:48]     = Conv_out[798];
    assign  image_1_65[47:32]     = Conv_out[770];
    assign  image_1_65[31:16]     = Conv_out[769];
    assign  image_1_65[15:0]      = Conv_out[768];

    assign  image_1_66[143:128]   = Conv_out[829];
    assign  image_1_66[127:112]   = Conv_out[828];
    assign  image_1_66[111:96]    = Conv_out[827];
    assign  image_1_66[95:80]     = Conv_out[799];
    assign  image_1_66[79:64]     = Conv_out[798];
    assign  image_1_66[63:48]     = Conv_out[797];
    assign  image_1_66[47:32]     = Conv_out[769];
    assign  image_1_66[31:16]     = Conv_out[768];
    assign  image_1_66[15:0]      = Conv_out[767];

    assign  image_1_67[143:128]   = Conv_out[828];
    assign  image_1_67[127:112]   = Conv_out[827];
    assign  image_1_67[111:96]    = Conv_out[826];
    assign  image_1_67[95:80]     = Conv_out[798];
    assign  image_1_67[79:64]     = Conv_out[797];
    assign  image_1_67[63:48]     = Conv_out[796];
    assign  image_1_67[47:32]     = Conv_out[768];
    assign  image_1_67[31:16]     = Conv_out[767];
    assign  image_1_67[15:0]      = Conv_out[766];

    assign  image_1_68[143:128]   = Conv_out[827];
    assign  image_1_68[127:112]   = Conv_out[826];
    assign  image_1_68[111:96]    = Conv_out[825];
    assign  image_1_68[95:80]     = Conv_out[797];
    assign  image_1_68[79:64]     = Conv_out[796];
    assign  image_1_68[63:48]     = Conv_out[795];
    assign  image_1_68[47:32]     = Conv_out[767];
    assign  image_1_68[31:16]     = Conv_out[766];
    assign  image_1_68[15:0]      = Conv_out[765];

    assign  image_1_69[143:128]   = Conv_out[826];
    assign  image_1_69[127:112]   = Conv_out[825];
    assign  image_1_69[111:96]    = Conv_out[824];
    assign  image_1_69[95:80]     = Conv_out[796];
    assign  image_1_69[79:64]     = Conv_out[795];
    assign  image_1_69[63:48]     = Conv_out[794];
    assign  image_1_69[47:32]     = Conv_out[766];
    assign  image_1_69[31:16]     = Conv_out[765];
    assign  image_1_69[15:0]      = Conv_out[764];

    assign  image_1_70[143:128]   = Conv_out[825];
    assign  image_1_70[127:112]   = Conv_out[824];
    assign  image_1_70[111:96]    = Conv_out[823];
    assign  image_1_70[95:80]     = Conv_out[795];
    assign  image_1_70[79:64]     = Conv_out[794];
    assign  image_1_70[63:48]     = Conv_out[793];
    assign  image_1_70[47:32]     = Conv_out[765];
    assign  image_1_70[31:16]     = Conv_out[764];
    assign  image_1_70[15:0]      = Conv_out[763];

    assign  image_1_71[143:128]   = Conv_out[824];
    assign  image_1_71[127:112]   = Conv_out[823];
    assign  image_1_71[111:96]    = Conv_out[822];
    assign  image_1_71[95:80]     = Conv_out[794];
    assign  image_1_71[79:64]     = Conv_out[793];
    assign  image_1_71[63:48]     = Conv_out[792];
    assign  image_1_71[47:32]     = Conv_out[764];
    assign  image_1_71[31:16]     = Conv_out[763];
    assign  image_1_71[15:0]      = Conv_out[762];

    assign  image_1_72[143:128]   = Conv_out[823];
    assign  image_1_72[127:112]   = Conv_out[822];
    assign  image_1_72[111:96]    = Conv_out[821];
    assign  image_1_72[95:80]     = Conv_out[793];
    assign  image_1_72[79:64]     = Conv_out[792];
    assign  image_1_72[63:48]     = Conv_out[791];
    assign  image_1_72[47:32]     = Conv_out[763];
    assign  image_1_72[31:16]     = Conv_out[762];
    assign  image_1_72[15:0]      = Conv_out[761];

    assign  image_1_73[143:128]   = Conv_out[822];
    assign  image_1_73[127:112]   = Conv_out[821];
    assign  image_1_73[111:96]    = Conv_out[820];
    assign  image_1_73[95:80]     = Conv_out[792];
    assign  image_1_73[79:64]     = Conv_out[791];
    assign  image_1_73[63:48]     = Conv_out[790];
    assign  image_1_73[47:32]     = Conv_out[762];
    assign  image_1_73[31:16]     = Conv_out[761];
    assign  image_1_73[15:0]      = Conv_out[760];

    assign  image_1_74[143:128]   = Conv_out[821];
    assign  image_1_74[127:112]   = Conv_out[820];
    assign  image_1_74[111:96]    = Conv_out[819];
    assign  image_1_74[95:80]     = Conv_out[791];
    assign  image_1_74[79:64]     = Conv_out[790];
    assign  image_1_74[63:48]     = Conv_out[789];
    assign  image_1_74[47:32]     = Conv_out[761];
    assign  image_1_74[31:16]     = Conv_out[760];
    assign  image_1_74[15:0]      = Conv_out[759];

    assign  image_1_75[143:128]   = Conv_out[820];
    assign  image_1_75[127:112]   = Conv_out[819];
    assign  image_1_75[111:96]    = Conv_out[818];
    assign  image_1_75[95:80]     = Conv_out[790];
    assign  image_1_75[79:64]     = Conv_out[789];
    assign  image_1_75[63:48]     = Conv_out[788];
    assign  image_1_75[47:32]     = Conv_out[760];
    assign  image_1_75[31:16]     = Conv_out[759];
    assign  image_1_75[15:0]      = Conv_out[758];

    assign  image_1_76[143:128]   = Conv_out[819];
    assign  image_1_76[127:112]   = Conv_out[818];
    assign  image_1_76[111:96]    = Conv_out[817];
    assign  image_1_76[95:80]     = Conv_out[789];
    assign  image_1_76[79:64]     = Conv_out[788];
    assign  image_1_76[63:48]     = Conv_out[787];
    assign  image_1_76[47:32]     = Conv_out[759];
    assign  image_1_76[31:16]     = Conv_out[758];
    assign  image_1_76[15:0]      = Conv_out[757];

    assign  image_1_77[143:128]   = Conv_out[818];
    assign  image_1_77[127:112]   = Conv_out[817];
    assign  image_1_77[111:96]    = Conv_out[816];
    assign  image_1_77[95:80]     = Conv_out[788];
    assign  image_1_77[79:64]     = Conv_out[787];
    assign  image_1_77[63:48]     = Conv_out[786];
    assign  image_1_77[47:32]     = Conv_out[758];
    assign  image_1_77[31:16]     = Conv_out[757];
    assign  image_1_77[15:0]      = Conv_out[756];

    assign  image_1_78[143:128]   = Conv_out[817];
    assign  image_1_78[127:112]   = Conv_out[816];
    assign  image_1_78[111:96]    = Conv_out[815];
    assign  image_1_78[95:80]     = Conv_out[787];
    assign  image_1_78[79:64]     = Conv_out[786];
    assign  image_1_78[63:48]     = Conv_out[785];
    assign  image_1_78[47:32]     = Conv_out[757];
    assign  image_1_78[31:16]     = Conv_out[756];
    assign  image_1_78[15:0]      = Conv_out[755];

    assign  image_1_79[143:128]   = Conv_out[816];
    assign  image_1_79[127:112]   = Conv_out[815];
    assign  image_1_79[111:96]    = Conv_out[814];
    assign  image_1_79[95:80]     = Conv_out[786];
    assign  image_1_79[79:64]     = Conv_out[785];
    assign  image_1_79[63:48]     = Conv_out[784];
    assign  image_1_79[47:32]     = Conv_out[756];
    assign  image_1_79[31:16]     = Conv_out[755];
    assign  image_1_79[15:0]      = Conv_out[754];

    assign  image_1_80[143:128]   = Conv_out[815];
    assign  image_1_80[127:112]   = Conv_out[814];
    assign  image_1_80[111:96]    = Conv_out[813];
    assign  image_1_80[95:80]     = Conv_out[785];
    assign  image_1_80[79:64]     = Conv_out[784];
    assign  image_1_80[63:48]     = Conv_out[783];
    assign  image_1_80[47:32]     = Conv_out[755];
    assign  image_1_80[31:16]     = Conv_out[754];
    assign  image_1_80[15:0]      = Conv_out[753];

    assign  image_1_81[143:128]   = Conv_out[814];
    assign  image_1_81[127:112]   = Conv_out[813];
    assign  image_1_81[111:96]    = Conv_out[812];
    assign  image_1_81[95:80]     = Conv_out[784];
    assign  image_1_81[79:64]     = Conv_out[783];
    assign  image_1_81[63:48]     = Conv_out[782];
    assign  image_1_81[47:32]     = Conv_out[754];
    assign  image_1_81[31:16]     = Conv_out[753];
    assign  image_1_81[15:0]      = Conv_out[752];

    assign  image_1_82[143:128]   = Conv_out[813];
    assign  image_1_82[127:112]   = Conv_out[812];
    assign  image_1_82[111:96]    = Conv_out[811];
    assign  image_1_82[95:80]     = Conv_out[783];
    assign  image_1_82[79:64]     = Conv_out[782];
    assign  image_1_82[63:48]     = Conv_out[781];
    assign  image_1_82[47:32]     = Conv_out[753];
    assign  image_1_82[31:16]     = Conv_out[752];
    assign  image_1_82[15:0]      = Conv_out[751];

    assign  image_1_83[143:128]   = Conv_out[812];
    assign  image_1_83[127:112]   = Conv_out[811];
    assign  image_1_83[111:96]    = Conv_out[810];
    assign  image_1_83[95:80]     = Conv_out[782];
    assign  image_1_83[79:64]     = Conv_out[781];
    assign  image_1_83[63:48]     = Conv_out[780];
    assign  image_1_83[47:32]     = Conv_out[752];
    assign  image_1_83[31:16]     = Conv_out[751];
    assign  image_1_83[15:0]      = Conv_out[750];

    assign  image_1_84[143:128]   = Conv_out[809];
    assign  image_1_84[127:112]   = Conv_out[808];
    assign  image_1_84[111:96]    = Conv_out[807];
    assign  image_1_84[95:80]     = Conv_out[779];
    assign  image_1_84[79:64]     = Conv_out[778];
    assign  image_1_84[63:48]     = Conv_out[777];
    assign  image_1_84[47:32]     = Conv_out[749];
    assign  image_1_84[31:16]     = Conv_out[748];
    assign  image_1_84[15:0]      = Conv_out[747];

    assign  image_1_85[143:128]   = Conv_out[808];
    assign  image_1_85[127:112]   = Conv_out[807];
    assign  image_1_85[111:96]    = Conv_out[806];
    assign  image_1_85[95:80]     = Conv_out[778];
    assign  image_1_85[79:64]     = Conv_out[777];
    assign  image_1_85[63:48]     = Conv_out[776];
    assign  image_1_85[47:32]     = Conv_out[748];
    assign  image_1_85[31:16]     = Conv_out[747];
    assign  image_1_85[15:0]      = Conv_out[746];

    assign  image_1_86[143:128]   = Conv_out[807];
    assign  image_1_86[127:112]   = Conv_out[806];
    assign  image_1_86[111:96]    = Conv_out[805];
    assign  image_1_86[95:80]     = Conv_out[777];
    assign  image_1_86[79:64]     = Conv_out[776];
    assign  image_1_86[63:48]     = Conv_out[775];
    assign  image_1_86[47:32]     = Conv_out[747];
    assign  image_1_86[31:16]     = Conv_out[746];
    assign  image_1_86[15:0]      = Conv_out[745];

    assign  image_1_87[143:128]   = Conv_out[806];
    assign  image_1_87[127:112]   = Conv_out[805];
    assign  image_1_87[111:96]    = Conv_out[804];
    assign  image_1_87[95:80]     = Conv_out[776];
    assign  image_1_87[79:64]     = Conv_out[775];
    assign  image_1_87[63:48]     = Conv_out[774];
    assign  image_1_87[47:32]     = Conv_out[746];
    assign  image_1_87[31:16]     = Conv_out[745];
    assign  image_1_87[15:0]      = Conv_out[744];

    assign  image_1_88[143:128]   = Conv_out[805];
    assign  image_1_88[127:112]   = Conv_out[804];
    assign  image_1_88[111:96]    = Conv_out[803];
    assign  image_1_88[95:80]     = Conv_out[775];
    assign  image_1_88[79:64]     = Conv_out[774];
    assign  image_1_88[63:48]     = Conv_out[773];
    assign  image_1_88[47:32]     = Conv_out[745];
    assign  image_1_88[31:16]     = Conv_out[744];
    assign  image_1_88[15:0]      = Conv_out[743];

    assign  image_1_89[143:128]   = Conv_out[804];
    assign  image_1_89[127:112]   = Conv_out[803];
    assign  image_1_89[111:96]    = Conv_out[802];
    assign  image_1_89[95:80]     = Conv_out[774];
    assign  image_1_89[79:64]     = Conv_out[773];
    assign  image_1_89[63:48]     = Conv_out[772];
    assign  image_1_89[47:32]     = Conv_out[744];
    assign  image_1_89[31:16]     = Conv_out[743];
    assign  image_1_89[15:0]      = Conv_out[742];

    assign  image_1_90[143:128]   = Conv_out[803];
    assign  image_1_90[127:112]   = Conv_out[802];
    assign  image_1_90[111:96]    = Conv_out[801];
    assign  image_1_90[95:80]     = Conv_out[773];
    assign  image_1_90[79:64]     = Conv_out[772];
    assign  image_1_90[63:48]     = Conv_out[771];
    assign  image_1_90[47:32]     = Conv_out[743];
    assign  image_1_90[31:16]     = Conv_out[742];
    assign  image_1_90[15:0]      = Conv_out[741];

    assign  image_1_91[143:128]   = Conv_out[802];
    assign  image_1_91[127:112]   = Conv_out[801];
    assign  image_1_91[111:96]    = Conv_out[800];
    assign  image_1_91[95:80]     = Conv_out[772];
    assign  image_1_91[79:64]     = Conv_out[771];
    assign  image_1_91[63:48]     = Conv_out[770];
    assign  image_1_91[47:32]     = Conv_out[742];
    assign  image_1_91[31:16]     = Conv_out[741];
    assign  image_1_91[15:0]      = Conv_out[740];

    assign  image_1_92[143:128]   = Conv_out[801];
    assign  image_1_92[127:112]   = Conv_out[800];
    assign  image_1_92[111:96]    = Conv_out[799];
    assign  image_1_92[95:80]     = Conv_out[771];
    assign  image_1_92[79:64]     = Conv_out[770];
    assign  image_1_92[63:48]     = Conv_out[769];
    assign  image_1_92[47:32]     = Conv_out[741];
    assign  image_1_92[31:16]     = Conv_out[740];
    assign  image_1_92[15:0]      = Conv_out[739];

    assign  image_1_93[143:128]   = Conv_out[800];
    assign  image_1_93[127:112]   = Conv_out[799];
    assign  image_1_93[111:96]    = Conv_out[798];
    assign  image_1_93[95:80]     = Conv_out[770];
    assign  image_1_93[79:64]     = Conv_out[769];
    assign  image_1_93[63:48]     = Conv_out[768];
    assign  image_1_93[47:32]     = Conv_out[740];
    assign  image_1_93[31:16]     = Conv_out[739];
    assign  image_1_93[15:0]      = Conv_out[738];

    assign  image_1_94[143:128]   = Conv_out[799];
    assign  image_1_94[127:112]   = Conv_out[798];
    assign  image_1_94[111:96]    = Conv_out[797];
    assign  image_1_94[95:80]     = Conv_out[769];
    assign  image_1_94[79:64]     = Conv_out[768];
    assign  image_1_94[63:48]     = Conv_out[767];
    assign  image_1_94[47:32]     = Conv_out[739];
    assign  image_1_94[31:16]     = Conv_out[738];
    assign  image_1_94[15:0]      = Conv_out[737];

    assign  image_1_95[143:128]   = Conv_out[798];
    assign  image_1_95[127:112]   = Conv_out[797];
    assign  image_1_95[111:96]    = Conv_out[796];
    assign  image_1_95[95:80]     = Conv_out[768];
    assign  image_1_95[79:64]     = Conv_out[767];
    assign  image_1_95[63:48]     = Conv_out[766];
    assign  image_1_95[47:32]     = Conv_out[738];
    assign  image_1_95[31:16]     = Conv_out[737];
    assign  image_1_95[15:0]      = Conv_out[736];

    assign  image_1_96[143:128]   = Conv_out[797];
    assign  image_1_96[127:112]   = Conv_out[796];
    assign  image_1_96[111:96]    = Conv_out[795];
    assign  image_1_96[95:80]     = Conv_out[767];
    assign  image_1_96[79:64]     = Conv_out[766];
    assign  image_1_96[63:48]     = Conv_out[765];
    assign  image_1_96[47:32]     = Conv_out[737];
    assign  image_1_96[31:16]     = Conv_out[736];
    assign  image_1_96[15:0]      = Conv_out[735];

    assign  image_1_97[143:128]   = Conv_out[796];
    assign  image_1_97[127:112]   = Conv_out[795];
    assign  image_1_97[111:96]    = Conv_out[794];
    assign  image_1_97[95:80]     = Conv_out[766];
    assign  image_1_97[79:64]     = Conv_out[765];
    assign  image_1_97[63:48]     = Conv_out[764];
    assign  image_1_97[47:32]     = Conv_out[736];
    assign  image_1_97[31:16]     = Conv_out[735];
    assign  image_1_97[15:0]      = Conv_out[734];

    assign  image_1_98[143:128]   = Conv_out[795];
    assign  image_1_98[127:112]   = Conv_out[794];
    assign  image_1_98[111:96]    = Conv_out[793];
    assign  image_1_98[95:80]     = Conv_out[765];
    assign  image_1_98[79:64]     = Conv_out[764];
    assign  image_1_98[63:48]     = Conv_out[763];
    assign  image_1_98[47:32]     = Conv_out[735];
    assign  image_1_98[31:16]     = Conv_out[734];
    assign  image_1_98[15:0]      = Conv_out[733];

    assign  image_1_99[143:128]   = Conv_out[794];
    assign  image_1_99[127:112]   = Conv_out[793];
    assign  image_1_99[111:96]    = Conv_out[792];
    assign  image_1_99[95:80]     = Conv_out[764];
    assign  image_1_99[79:64]     = Conv_out[763];
    assign  image_1_99[63:48]     = Conv_out[762];
    assign  image_1_99[47:32]     = Conv_out[734];
    assign  image_1_99[31:16]     = Conv_out[733];
    assign  image_1_99[15:0]      = Conv_out[732];

    assign  image_1_100[143:128]   = Conv_out[793];
    assign  image_1_100[127:112]   = Conv_out[792];
    assign  image_1_100[111:96]    = Conv_out[791];
    assign  image_1_100[95:80]     = Conv_out[763];
    assign  image_1_100[79:64]     = Conv_out[762];
    assign  image_1_100[63:48]     = Conv_out[761];
    assign  image_1_100[47:32]     = Conv_out[733];
    assign  image_1_100[31:16]     = Conv_out[732];
    assign  image_1_100[15:0]      = Conv_out[731];

    assign  image_1_101[143:128]   = Conv_out[792];
    assign  image_1_101[127:112]   = Conv_out[791];
    assign  image_1_101[111:96]    = Conv_out[790];
    assign  image_1_101[95:80]     = Conv_out[762];
    assign  image_1_101[79:64]     = Conv_out[761];
    assign  image_1_101[63:48]     = Conv_out[760];
    assign  image_1_101[47:32]     = Conv_out[732];
    assign  image_1_101[31:16]     = Conv_out[731];
    assign  image_1_101[15:0]      = Conv_out[730];

    assign  image_1_102[143:128]   = Conv_out[791];
    assign  image_1_102[127:112]   = Conv_out[790];
    assign  image_1_102[111:96]    = Conv_out[789];
    assign  image_1_102[95:80]     = Conv_out[761];
    assign  image_1_102[79:64]     = Conv_out[760];
    assign  image_1_102[63:48]     = Conv_out[759];
    assign  image_1_102[47:32]     = Conv_out[731];
    assign  image_1_102[31:16]     = Conv_out[730];
    assign  image_1_102[15:0]      = Conv_out[729];

    assign  image_1_103[143:128]   = Conv_out[790];
    assign  image_1_103[127:112]   = Conv_out[789];
    assign  image_1_103[111:96]    = Conv_out[788];
    assign  image_1_103[95:80]     = Conv_out[760];
    assign  image_1_103[79:64]     = Conv_out[759];
    assign  image_1_103[63:48]     = Conv_out[758];
    assign  image_1_103[47:32]     = Conv_out[730];
    assign  image_1_103[31:16]     = Conv_out[729];
    assign  image_1_103[15:0]      = Conv_out[728];

    assign  image_1_104[143:128]   = Conv_out[789];
    assign  image_1_104[127:112]   = Conv_out[788];
    assign  image_1_104[111:96]    = Conv_out[787];
    assign  image_1_104[95:80]     = Conv_out[759];
    assign  image_1_104[79:64]     = Conv_out[758];
    assign  image_1_104[63:48]     = Conv_out[757];
    assign  image_1_104[47:32]     = Conv_out[729];
    assign  image_1_104[31:16]     = Conv_out[728];
    assign  image_1_104[15:0]      = Conv_out[727];

    assign  image_1_105[143:128]   = Conv_out[788];
    assign  image_1_105[127:112]   = Conv_out[787];
    assign  image_1_105[111:96]    = Conv_out[786];
    assign  image_1_105[95:80]     = Conv_out[758];
    assign  image_1_105[79:64]     = Conv_out[757];
    assign  image_1_105[63:48]     = Conv_out[756];
    assign  image_1_105[47:32]     = Conv_out[728];
    assign  image_1_105[31:16]     = Conv_out[727];
    assign  image_1_105[15:0]      = Conv_out[726];

    assign  image_1_106[143:128]   = Conv_out[787];
    assign  image_1_106[127:112]   = Conv_out[786];
    assign  image_1_106[111:96]    = Conv_out[785];
    assign  image_1_106[95:80]     = Conv_out[757];
    assign  image_1_106[79:64]     = Conv_out[756];
    assign  image_1_106[63:48]     = Conv_out[755];
    assign  image_1_106[47:32]     = Conv_out[727];
    assign  image_1_106[31:16]     = Conv_out[726];
    assign  image_1_106[15:0]      = Conv_out[725];

    assign  image_1_107[143:128]   = Conv_out[786];
    assign  image_1_107[127:112]   = Conv_out[785];
    assign  image_1_107[111:96]    = Conv_out[784];
    assign  image_1_107[95:80]     = Conv_out[756];
    assign  image_1_107[79:64]     = Conv_out[755];
    assign  image_1_107[63:48]     = Conv_out[754];
    assign  image_1_107[47:32]     = Conv_out[726];
    assign  image_1_107[31:16]     = Conv_out[725];
    assign  image_1_107[15:0]      = Conv_out[724];

    assign  image_1_108[143:128]   = Conv_out[785];
    assign  image_1_108[127:112]   = Conv_out[784];
    assign  image_1_108[111:96]    = Conv_out[783];
    assign  image_1_108[95:80]     = Conv_out[755];
    assign  image_1_108[79:64]     = Conv_out[754];
    assign  image_1_108[63:48]     = Conv_out[753];
    assign  image_1_108[47:32]     = Conv_out[725];
    assign  image_1_108[31:16]     = Conv_out[724];
    assign  image_1_108[15:0]      = Conv_out[723];

    assign  image_1_109[143:128]   = Conv_out[784];
    assign  image_1_109[127:112]   = Conv_out[783];
    assign  image_1_109[111:96]    = Conv_out[782];
    assign  image_1_109[95:80]     = Conv_out[754];
    assign  image_1_109[79:64]     = Conv_out[753];
    assign  image_1_109[63:48]     = Conv_out[752];
    assign  image_1_109[47:32]     = Conv_out[724];
    assign  image_1_109[31:16]     = Conv_out[723];
    assign  image_1_109[15:0]      = Conv_out[722];

    assign  image_1_110[143:128]   = Conv_out[783];
    assign  image_1_110[127:112]   = Conv_out[782];
    assign  image_1_110[111:96]    = Conv_out[781];
    assign  image_1_110[95:80]     = Conv_out[753];
    assign  image_1_110[79:64]     = Conv_out[752];
    assign  image_1_110[63:48]     = Conv_out[751];
    assign  image_1_110[47:32]     = Conv_out[723];
    assign  image_1_110[31:16]     = Conv_out[722];
    assign  image_1_110[15:0]      = Conv_out[721];

    assign  image_1_111[143:128]   = Conv_out[782];
    assign  image_1_111[127:112]   = Conv_out[781];
    assign  image_1_111[111:96]    = Conv_out[780];
    assign  image_1_111[95:80]     = Conv_out[752];
    assign  image_1_111[79:64]     = Conv_out[751];
    assign  image_1_111[63:48]     = Conv_out[750];
    assign  image_1_111[47:32]     = Conv_out[722];
    assign  image_1_111[31:16]     = Conv_out[721];
    assign  image_1_111[15:0]      = Conv_out[720];

    assign  image_1_112[143:128]   = Conv_out[779];
    assign  image_1_112[127:112]   = Conv_out[778];
    assign  image_1_112[111:96]    = Conv_out[777];
    assign  image_1_112[95:80]     = Conv_out[749];
    assign  image_1_112[79:64]     = Conv_out[748];
    assign  image_1_112[63:48]     = Conv_out[747];
    assign  image_1_112[47:32]     = Conv_out[719];
    assign  image_1_112[31:16]     = Conv_out[718];
    assign  image_1_112[15:0]      = Conv_out[717];

    assign  image_1_113[143:128]   = Conv_out[778];
    assign  image_1_113[127:112]   = Conv_out[777];
    assign  image_1_113[111:96]    = Conv_out[776];
    assign  image_1_113[95:80]     = Conv_out[748];
    assign  image_1_113[79:64]     = Conv_out[747];
    assign  image_1_113[63:48]     = Conv_out[746];
    assign  image_1_113[47:32]     = Conv_out[718];
    assign  image_1_113[31:16]     = Conv_out[717];
    assign  image_1_113[15:0]      = Conv_out[716];

    assign  image_1_114[143:128]   = Conv_out[777];
    assign  image_1_114[127:112]   = Conv_out[776];
    assign  image_1_114[111:96]    = Conv_out[775];
    assign  image_1_114[95:80]     = Conv_out[747];
    assign  image_1_114[79:64]     = Conv_out[746];
    assign  image_1_114[63:48]     = Conv_out[745];
    assign  image_1_114[47:32]     = Conv_out[717];
    assign  image_1_114[31:16]     = Conv_out[716];
    assign  image_1_114[15:0]      = Conv_out[715];

    assign  image_1_115[143:128]   = Conv_out[776];
    assign  image_1_115[127:112]   = Conv_out[775];
    assign  image_1_115[111:96]    = Conv_out[774];
    assign  image_1_115[95:80]     = Conv_out[746];
    assign  image_1_115[79:64]     = Conv_out[745];
    assign  image_1_115[63:48]     = Conv_out[744];
    assign  image_1_115[47:32]     = Conv_out[716];
    assign  image_1_115[31:16]     = Conv_out[715];
    assign  image_1_115[15:0]      = Conv_out[714];

    assign  image_1_116[143:128]   = Conv_out[775];
    assign  image_1_116[127:112]   = Conv_out[774];
    assign  image_1_116[111:96]    = Conv_out[773];
    assign  image_1_116[95:80]     = Conv_out[745];
    assign  image_1_116[79:64]     = Conv_out[744];
    assign  image_1_116[63:48]     = Conv_out[743];
    assign  image_1_116[47:32]     = Conv_out[715];
    assign  image_1_116[31:16]     = Conv_out[714];
    assign  image_1_116[15:0]      = Conv_out[713];

    assign  image_1_117[143:128]   = Conv_out[774];
    assign  image_1_117[127:112]   = Conv_out[773];
    assign  image_1_117[111:96]    = Conv_out[772];
    assign  image_1_117[95:80]     = Conv_out[744];
    assign  image_1_117[79:64]     = Conv_out[743];
    assign  image_1_117[63:48]     = Conv_out[742];
    assign  image_1_117[47:32]     = Conv_out[714];
    assign  image_1_117[31:16]     = Conv_out[713];
    assign  image_1_117[15:0]      = Conv_out[712];

    assign  image_1_118[143:128]   = Conv_out[773];
    assign  image_1_118[127:112]   = Conv_out[772];
    assign  image_1_118[111:96]    = Conv_out[771];
    assign  image_1_118[95:80]     = Conv_out[743];
    assign  image_1_118[79:64]     = Conv_out[742];
    assign  image_1_118[63:48]     = Conv_out[741];
    assign  image_1_118[47:32]     = Conv_out[713];
    assign  image_1_118[31:16]     = Conv_out[712];
    assign  image_1_118[15:0]      = Conv_out[711];

    assign  image_1_119[143:128]   = Conv_out[772];
    assign  image_1_119[127:112]   = Conv_out[771];
    assign  image_1_119[111:96]    = Conv_out[770];
    assign  image_1_119[95:80]     = Conv_out[742];
    assign  image_1_119[79:64]     = Conv_out[741];
    assign  image_1_119[63:48]     = Conv_out[740];
    assign  image_1_119[47:32]     = Conv_out[712];
    assign  image_1_119[31:16]     = Conv_out[711];
    assign  image_1_119[15:0]      = Conv_out[710];

    assign  image_1_120[143:128]   = Conv_out[771];
    assign  image_1_120[127:112]   = Conv_out[770];
    assign  image_1_120[111:96]    = Conv_out[769];
    assign  image_1_120[95:80]     = Conv_out[741];
    assign  image_1_120[79:64]     = Conv_out[740];
    assign  image_1_120[63:48]     = Conv_out[739];
    assign  image_1_120[47:32]     = Conv_out[711];
    assign  image_1_120[31:16]     = Conv_out[710];
    assign  image_1_120[15:0]      = Conv_out[709];

    assign  image_1_121[143:128]   = Conv_out[770];
    assign  image_1_121[127:112]   = Conv_out[769];
    assign  image_1_121[111:96]    = Conv_out[768];
    assign  image_1_121[95:80]     = Conv_out[740];
    assign  image_1_121[79:64]     = Conv_out[739];
    assign  image_1_121[63:48]     = Conv_out[738];
    assign  image_1_121[47:32]     = Conv_out[710];
    assign  image_1_121[31:16]     = Conv_out[709];
    assign  image_1_121[15:0]      = Conv_out[708];

    assign  image_1_122[143:128]   = Conv_out[769];
    assign  image_1_122[127:112]   = Conv_out[768];
    assign  image_1_122[111:96]    = Conv_out[767];
    assign  image_1_122[95:80]     = Conv_out[739];
    assign  image_1_122[79:64]     = Conv_out[738];
    assign  image_1_122[63:48]     = Conv_out[737];
    assign  image_1_122[47:32]     = Conv_out[709];
    assign  image_1_122[31:16]     = Conv_out[708];
    assign  image_1_122[15:0]      = Conv_out[707];

    assign  image_1_123[143:128]   = Conv_out[768];
    assign  image_1_123[127:112]   = Conv_out[767];
    assign  image_1_123[111:96]    = Conv_out[766];
    assign  image_1_123[95:80]     = Conv_out[738];
    assign  image_1_123[79:64]     = Conv_out[737];
    assign  image_1_123[63:48]     = Conv_out[736];
    assign  image_1_123[47:32]     = Conv_out[708];
    assign  image_1_123[31:16]     = Conv_out[707];
    assign  image_1_123[15:0]      = Conv_out[706];

    assign  image_1_124[143:128]   = Conv_out[767];
    assign  image_1_124[127:112]   = Conv_out[766];
    assign  image_1_124[111:96]    = Conv_out[765];
    assign  image_1_124[95:80]     = Conv_out[737];
    assign  image_1_124[79:64]     = Conv_out[736];
    assign  image_1_124[63:48]     = Conv_out[735];
    assign  image_1_124[47:32]     = Conv_out[707];
    assign  image_1_124[31:16]     = Conv_out[706];
    assign  image_1_124[15:0]      = Conv_out[705];

    assign  image_1_125[143:128]   = Conv_out[766];
    assign  image_1_125[127:112]   = Conv_out[765];
    assign  image_1_125[111:96]    = Conv_out[764];
    assign  image_1_125[95:80]     = Conv_out[736];
    assign  image_1_125[79:64]     = Conv_out[735];
    assign  image_1_125[63:48]     = Conv_out[734];
    assign  image_1_125[47:32]     = Conv_out[706];
    assign  image_1_125[31:16]     = Conv_out[705];
    assign  image_1_125[15:0]      = Conv_out[704];

    assign  image_1_126[143:128]   = Conv_out[765];
    assign  image_1_126[127:112]   = Conv_out[764];
    assign  image_1_126[111:96]    = Conv_out[763];
    assign  image_1_126[95:80]     = Conv_out[735];
    assign  image_1_126[79:64]     = Conv_out[734];
    assign  image_1_126[63:48]     = Conv_out[733];
    assign  image_1_126[47:32]     = Conv_out[705];
    assign  image_1_126[31:16]     = Conv_out[704];
    assign  image_1_126[15:0]      = Conv_out[703];

    assign  image_1_127[143:128]   = Conv_out[764];
    assign  image_1_127[127:112]   = Conv_out[763];
    assign  image_1_127[111:96]    = Conv_out[762];
    assign  image_1_127[95:80]     = Conv_out[734];
    assign  image_1_127[79:64]     = Conv_out[733];
    assign  image_1_127[63:48]     = Conv_out[732];
    assign  image_1_127[47:32]     = Conv_out[704];
    assign  image_1_127[31:16]     = Conv_out[703];
    assign  image_1_127[15:0]      = Conv_out[702];

    assign  image_1_128[143:128]   = Conv_out[763];
    assign  image_1_128[127:112]   = Conv_out[762];
    assign  image_1_128[111:96]    = Conv_out[761];
    assign  image_1_128[95:80]     = Conv_out[733];
    assign  image_1_128[79:64]     = Conv_out[732];
    assign  image_1_128[63:48]     = Conv_out[731];
    assign  image_1_128[47:32]     = Conv_out[703];
    assign  image_1_128[31:16]     = Conv_out[702];
    assign  image_1_128[15:0]      = Conv_out[701];

    assign  image_1_129[143:128]   = Conv_out[762];
    assign  image_1_129[127:112]   = Conv_out[761];
    assign  image_1_129[111:96]    = Conv_out[760];
    assign  image_1_129[95:80]     = Conv_out[732];
    assign  image_1_129[79:64]     = Conv_out[731];
    assign  image_1_129[63:48]     = Conv_out[730];
    assign  image_1_129[47:32]     = Conv_out[702];
    assign  image_1_129[31:16]     = Conv_out[701];
    assign  image_1_129[15:0]      = Conv_out[700];

    assign  image_1_130[143:128]   = Conv_out[761];
    assign  image_1_130[127:112]   = Conv_out[760];
    assign  image_1_130[111:96]    = Conv_out[759];
    assign  image_1_130[95:80]     = Conv_out[731];
    assign  image_1_130[79:64]     = Conv_out[730];
    assign  image_1_130[63:48]     = Conv_out[729];
    assign  image_1_130[47:32]     = Conv_out[701];
    assign  image_1_130[31:16]     = Conv_out[700];
    assign  image_1_130[15:0]      = Conv_out[699];

    assign  image_1_131[143:128]   = Conv_out[760];
    assign  image_1_131[127:112]   = Conv_out[759];
    assign  image_1_131[111:96]    = Conv_out[758];
    assign  image_1_131[95:80]     = Conv_out[730];
    assign  image_1_131[79:64]     = Conv_out[729];
    assign  image_1_131[63:48]     = Conv_out[728];
    assign  image_1_131[47:32]     = Conv_out[700];
    assign  image_1_131[31:16]     = Conv_out[699];
    assign  image_1_131[15:0]      = Conv_out[698];

    assign  image_1_132[143:128]   = Conv_out[759];
    assign  image_1_132[127:112]   = Conv_out[758];
    assign  image_1_132[111:96]    = Conv_out[757];
    assign  image_1_132[95:80]     = Conv_out[729];
    assign  image_1_132[79:64]     = Conv_out[728];
    assign  image_1_132[63:48]     = Conv_out[727];
    assign  image_1_132[47:32]     = Conv_out[699];
    assign  image_1_132[31:16]     = Conv_out[698];
    assign  image_1_132[15:0]      = Conv_out[697];

    assign  image_1_133[143:128]   = Conv_out[758];
    assign  image_1_133[127:112]   = Conv_out[757];
    assign  image_1_133[111:96]    = Conv_out[756];
    assign  image_1_133[95:80]     = Conv_out[728];
    assign  image_1_133[79:64]     = Conv_out[727];
    assign  image_1_133[63:48]     = Conv_out[726];
    assign  image_1_133[47:32]     = Conv_out[698];
    assign  image_1_133[31:16]     = Conv_out[697];
    assign  image_1_133[15:0]      = Conv_out[696];

    assign  image_1_134[143:128]   = Conv_out[757];
    assign  image_1_134[127:112]   = Conv_out[756];
    assign  image_1_134[111:96]    = Conv_out[755];
    assign  image_1_134[95:80]     = Conv_out[727];
    assign  image_1_134[79:64]     = Conv_out[726];
    assign  image_1_134[63:48]     = Conv_out[725];
    assign  image_1_134[47:32]     = Conv_out[697];
    assign  image_1_134[31:16]     = Conv_out[696];
    assign  image_1_134[15:0]      = Conv_out[695];

    assign  image_1_135[143:128]   = Conv_out[756];
    assign  image_1_135[127:112]   = Conv_out[755];
    assign  image_1_135[111:96]    = Conv_out[754];
    assign  image_1_135[95:80]     = Conv_out[726];
    assign  image_1_135[79:64]     = Conv_out[725];
    assign  image_1_135[63:48]     = Conv_out[724];
    assign  image_1_135[47:32]     = Conv_out[696];
    assign  image_1_135[31:16]     = Conv_out[695];
    assign  image_1_135[15:0]      = Conv_out[694];

    assign  image_1_136[143:128]   = Conv_out[755];
    assign  image_1_136[127:112]   = Conv_out[754];
    assign  image_1_136[111:96]    = Conv_out[753];
    assign  image_1_136[95:80]     = Conv_out[725];
    assign  image_1_136[79:64]     = Conv_out[724];
    assign  image_1_136[63:48]     = Conv_out[723];
    assign  image_1_136[47:32]     = Conv_out[695];
    assign  image_1_136[31:16]     = Conv_out[694];
    assign  image_1_136[15:0]      = Conv_out[693];

    assign  image_1_137[143:128]   = Conv_out[754];
    assign  image_1_137[127:112]   = Conv_out[753];
    assign  image_1_137[111:96]    = Conv_out[752];
    assign  image_1_137[95:80]     = Conv_out[724];
    assign  image_1_137[79:64]     = Conv_out[723];
    assign  image_1_137[63:48]     = Conv_out[722];
    assign  image_1_137[47:32]     = Conv_out[694];
    assign  image_1_137[31:16]     = Conv_out[693];
    assign  image_1_137[15:0]      = Conv_out[692];

    assign  image_1_138[143:128]   = Conv_out[753];
    assign  image_1_138[127:112]   = Conv_out[752];
    assign  image_1_138[111:96]    = Conv_out[751];
    assign  image_1_138[95:80]     = Conv_out[723];
    assign  image_1_138[79:64]     = Conv_out[722];
    assign  image_1_138[63:48]     = Conv_out[721];
    assign  image_1_138[47:32]     = Conv_out[693];
    assign  image_1_138[31:16]     = Conv_out[692];
    assign  image_1_138[15:0]      = Conv_out[691];

    assign  image_1_139[143:128]   = Conv_out[752];
    assign  image_1_139[127:112]   = Conv_out[751];
    assign  image_1_139[111:96]    = Conv_out[750];
    assign  image_1_139[95:80]     = Conv_out[722];
    assign  image_1_139[79:64]     = Conv_out[721];
    assign  image_1_139[63:48]     = Conv_out[720];
    assign  image_1_139[47:32]     = Conv_out[692];
    assign  image_1_139[31:16]     = Conv_out[691];
    assign  image_1_139[15:0]      = Conv_out[690];

    assign  image_1_140[143:128]   = Conv_out[749];
    assign  image_1_140[127:112]   = Conv_out[748];
    assign  image_1_140[111:96]    = Conv_out[747];
    assign  image_1_140[95:80]     = Conv_out[719];
    assign  image_1_140[79:64]     = Conv_out[718];
    assign  image_1_140[63:48]     = Conv_out[717];
    assign  image_1_140[47:32]     = Conv_out[689];
    assign  image_1_140[31:16]     = Conv_out[688];
    assign  image_1_140[15:0]      = Conv_out[687];

    assign  image_1_141[143:128]   = Conv_out[748];
    assign  image_1_141[127:112]   = Conv_out[747];
    assign  image_1_141[111:96]    = Conv_out[746];
    assign  image_1_141[95:80]     = Conv_out[718];
    assign  image_1_141[79:64]     = Conv_out[717];
    assign  image_1_141[63:48]     = Conv_out[716];
    assign  image_1_141[47:32]     = Conv_out[688];
    assign  image_1_141[31:16]     = Conv_out[687];
    assign  image_1_141[15:0]      = Conv_out[686];

    assign  image_1_142[143:128]   = Conv_out[747];
    assign  image_1_142[127:112]   = Conv_out[746];
    assign  image_1_142[111:96]    = Conv_out[745];
    assign  image_1_142[95:80]     = Conv_out[717];
    assign  image_1_142[79:64]     = Conv_out[716];
    assign  image_1_142[63:48]     = Conv_out[715];
    assign  image_1_142[47:32]     = Conv_out[687];
    assign  image_1_142[31:16]     = Conv_out[686];
    assign  image_1_142[15:0]      = Conv_out[685];

    assign  image_1_143[143:128]   = Conv_out[746];
    assign  image_1_143[127:112]   = Conv_out[745];
    assign  image_1_143[111:96]    = Conv_out[744];
    assign  image_1_143[95:80]     = Conv_out[716];
    assign  image_1_143[79:64]     = Conv_out[715];
    assign  image_1_143[63:48]     = Conv_out[714];
    assign  image_1_143[47:32]     = Conv_out[686];
    assign  image_1_143[31:16]     = Conv_out[685];
    assign  image_1_143[15:0]      = Conv_out[684];

    assign  image_1_144[143:128]   = Conv_out[745];
    assign  image_1_144[127:112]   = Conv_out[744];
    assign  image_1_144[111:96]    = Conv_out[743];
    assign  image_1_144[95:80]     = Conv_out[715];
    assign  image_1_144[79:64]     = Conv_out[714];
    assign  image_1_144[63:48]     = Conv_out[713];
    assign  image_1_144[47:32]     = Conv_out[685];
    assign  image_1_144[31:16]     = Conv_out[684];
    assign  image_1_144[15:0]      = Conv_out[683];

    assign  image_1_145[143:128]   = Conv_out[744];
    assign  image_1_145[127:112]   = Conv_out[743];
    assign  image_1_145[111:96]    = Conv_out[742];
    assign  image_1_145[95:80]     = Conv_out[714];
    assign  image_1_145[79:64]     = Conv_out[713];
    assign  image_1_145[63:48]     = Conv_out[712];
    assign  image_1_145[47:32]     = Conv_out[684];
    assign  image_1_145[31:16]     = Conv_out[683];
    assign  image_1_145[15:0]      = Conv_out[682];

    assign  image_1_146[143:128]   = Conv_out[743];
    assign  image_1_146[127:112]   = Conv_out[742];
    assign  image_1_146[111:96]    = Conv_out[741];
    assign  image_1_146[95:80]     = Conv_out[713];
    assign  image_1_146[79:64]     = Conv_out[712];
    assign  image_1_146[63:48]     = Conv_out[711];
    assign  image_1_146[47:32]     = Conv_out[683];
    assign  image_1_146[31:16]     = Conv_out[682];
    assign  image_1_146[15:0]      = Conv_out[681];

    assign  image_1_147[143:128]   = Conv_out[742];
    assign  image_1_147[127:112]   = Conv_out[741];
    assign  image_1_147[111:96]    = Conv_out[740];
    assign  image_1_147[95:80]     = Conv_out[712];
    assign  image_1_147[79:64]     = Conv_out[711];
    assign  image_1_147[63:48]     = Conv_out[710];
    assign  image_1_147[47:32]     = Conv_out[682];
    assign  image_1_147[31:16]     = Conv_out[681];
    assign  image_1_147[15:0]      = Conv_out[680];

    assign  image_1_148[143:128]   = Conv_out[741];
    assign  image_1_148[127:112]   = Conv_out[740];
    assign  image_1_148[111:96]    = Conv_out[739];
    assign  image_1_148[95:80]     = Conv_out[711];
    assign  image_1_148[79:64]     = Conv_out[710];
    assign  image_1_148[63:48]     = Conv_out[709];
    assign  image_1_148[47:32]     = Conv_out[681];
    assign  image_1_148[31:16]     = Conv_out[680];
    assign  image_1_148[15:0]      = Conv_out[679];

    assign  image_1_149[143:128]   = Conv_out[740];
    assign  image_1_149[127:112]   = Conv_out[739];
    assign  image_1_149[111:96]    = Conv_out[738];
    assign  image_1_149[95:80]     = Conv_out[710];
    assign  image_1_149[79:64]     = Conv_out[709];
    assign  image_1_149[63:48]     = Conv_out[708];
    assign  image_1_149[47:32]     = Conv_out[680];
    assign  image_1_149[31:16]     = Conv_out[679];
    assign  image_1_149[15:0]      = Conv_out[678];

    assign  image_1_150[143:128]   = Conv_out[739];
    assign  image_1_150[127:112]   = Conv_out[738];
    assign  image_1_150[111:96]    = Conv_out[737];
    assign  image_1_150[95:80]     = Conv_out[709];
    assign  image_1_150[79:64]     = Conv_out[708];
    assign  image_1_150[63:48]     = Conv_out[707];
    assign  image_1_150[47:32]     = Conv_out[679];
    assign  image_1_150[31:16]     = Conv_out[678];
    assign  image_1_150[15:0]      = Conv_out[677];

    assign  image_1_151[143:128]   = Conv_out[738];
    assign  image_1_151[127:112]   = Conv_out[737];
    assign  image_1_151[111:96]    = Conv_out[736];
    assign  image_1_151[95:80]     = Conv_out[708];
    assign  image_1_151[79:64]     = Conv_out[707];
    assign  image_1_151[63:48]     = Conv_out[706];
    assign  image_1_151[47:32]     = Conv_out[678];
    assign  image_1_151[31:16]     = Conv_out[677];
    assign  image_1_151[15:0]      = Conv_out[676];

    assign  image_1_152[143:128]   = Conv_out[737];
    assign  image_1_152[127:112]   = Conv_out[736];
    assign  image_1_152[111:96]    = Conv_out[735];
    assign  image_1_152[95:80]     = Conv_out[707];
    assign  image_1_152[79:64]     = Conv_out[706];
    assign  image_1_152[63:48]     = Conv_out[705];
    assign  image_1_152[47:32]     = Conv_out[677];
    assign  image_1_152[31:16]     = Conv_out[676];
    assign  image_1_152[15:0]      = Conv_out[675];

    assign  image_1_153[143:128]   = Conv_out[736];
    assign  image_1_153[127:112]   = Conv_out[735];
    assign  image_1_153[111:96]    = Conv_out[734];
    assign  image_1_153[95:80]     = Conv_out[706];
    assign  image_1_153[79:64]     = Conv_out[705];
    assign  image_1_153[63:48]     = Conv_out[704];
    assign  image_1_153[47:32]     = Conv_out[676];
    assign  image_1_153[31:16]     = Conv_out[675];
    assign  image_1_153[15:0]      = Conv_out[674];

    assign  image_1_154[143:128]   = Conv_out[735];
    assign  image_1_154[127:112]   = Conv_out[734];
    assign  image_1_154[111:96]    = Conv_out[733];
    assign  image_1_154[95:80]     = Conv_out[705];
    assign  image_1_154[79:64]     = Conv_out[704];
    assign  image_1_154[63:48]     = Conv_out[703];
    assign  image_1_154[47:32]     = Conv_out[675];
    assign  image_1_154[31:16]     = Conv_out[674];
    assign  image_1_154[15:0]      = Conv_out[673];

    assign  image_1_155[143:128]   = Conv_out[734];
    assign  image_1_155[127:112]   = Conv_out[733];
    assign  image_1_155[111:96]    = Conv_out[732];
    assign  image_1_155[95:80]     = Conv_out[704];
    assign  image_1_155[79:64]     = Conv_out[703];
    assign  image_1_155[63:48]     = Conv_out[702];
    assign  image_1_155[47:32]     = Conv_out[674];
    assign  image_1_155[31:16]     = Conv_out[673];
    assign  image_1_155[15:0]      = Conv_out[672];

    assign  image_1_156[143:128]   = Conv_out[733];
    assign  image_1_156[127:112]   = Conv_out[732];
    assign  image_1_156[111:96]    = Conv_out[731];
    assign  image_1_156[95:80]     = Conv_out[703];
    assign  image_1_156[79:64]     = Conv_out[702];
    assign  image_1_156[63:48]     = Conv_out[701];
    assign  image_1_156[47:32]     = Conv_out[673];
    assign  image_1_156[31:16]     = Conv_out[672];
    assign  image_1_156[15:0]      = Conv_out[671];

    assign  image_1_157[143:128]   = Conv_out[732];
    assign  image_1_157[127:112]   = Conv_out[731];
    assign  image_1_157[111:96]    = Conv_out[730];
    assign  image_1_157[95:80]     = Conv_out[702];
    assign  image_1_157[79:64]     = Conv_out[701];
    assign  image_1_157[63:48]     = Conv_out[700];
    assign  image_1_157[47:32]     = Conv_out[672];
    assign  image_1_157[31:16]     = Conv_out[671];
    assign  image_1_157[15:0]      = Conv_out[670];

    assign  image_1_158[143:128]   = Conv_out[731];
    assign  image_1_158[127:112]   = Conv_out[730];
    assign  image_1_158[111:96]    = Conv_out[729];
    assign  image_1_158[95:80]     = Conv_out[701];
    assign  image_1_158[79:64]     = Conv_out[700];
    assign  image_1_158[63:48]     = Conv_out[699];
    assign  image_1_158[47:32]     = Conv_out[671];
    assign  image_1_158[31:16]     = Conv_out[670];
    assign  image_1_158[15:0]      = Conv_out[669];

    assign  image_1_159[143:128]   = Conv_out[730];
    assign  image_1_159[127:112]   = Conv_out[729];
    assign  image_1_159[111:96]    = Conv_out[728];
    assign  image_1_159[95:80]     = Conv_out[700];
    assign  image_1_159[79:64]     = Conv_out[699];
    assign  image_1_159[63:48]     = Conv_out[698];
    assign  image_1_159[47:32]     = Conv_out[670];
    assign  image_1_159[31:16]     = Conv_out[669];
    assign  image_1_159[15:0]      = Conv_out[668];

    assign  image_1_160[143:128]   = Conv_out[729];
    assign  image_1_160[127:112]   = Conv_out[728];
    assign  image_1_160[111:96]    = Conv_out[727];
    assign  image_1_160[95:80]     = Conv_out[699];
    assign  image_1_160[79:64]     = Conv_out[698];
    assign  image_1_160[63:48]     = Conv_out[697];
    assign  image_1_160[47:32]     = Conv_out[669];
    assign  image_1_160[31:16]     = Conv_out[668];
    assign  image_1_160[15:0]      = Conv_out[667];

    assign  image_1_161[143:128]   = Conv_out[728];
    assign  image_1_161[127:112]   = Conv_out[727];
    assign  image_1_161[111:96]    = Conv_out[726];
    assign  image_1_161[95:80]     = Conv_out[698];
    assign  image_1_161[79:64]     = Conv_out[697];
    assign  image_1_161[63:48]     = Conv_out[696];
    assign  image_1_161[47:32]     = Conv_out[668];
    assign  image_1_161[31:16]     = Conv_out[667];
    assign  image_1_161[15:0]      = Conv_out[666];

    assign  image_1_162[143:128]   = Conv_out[727];
    assign  image_1_162[127:112]   = Conv_out[726];
    assign  image_1_162[111:96]    = Conv_out[725];
    assign  image_1_162[95:80]     = Conv_out[697];
    assign  image_1_162[79:64]     = Conv_out[696];
    assign  image_1_162[63:48]     = Conv_out[695];
    assign  image_1_162[47:32]     = Conv_out[667];
    assign  image_1_162[31:16]     = Conv_out[666];
    assign  image_1_162[15:0]      = Conv_out[665];

    assign  image_1_163[143:128]   = Conv_out[726];
    assign  image_1_163[127:112]   = Conv_out[725];
    assign  image_1_163[111:96]    = Conv_out[724];
    assign  image_1_163[95:80]     = Conv_out[696];
    assign  image_1_163[79:64]     = Conv_out[695];
    assign  image_1_163[63:48]     = Conv_out[694];
    assign  image_1_163[47:32]     = Conv_out[666];
    assign  image_1_163[31:16]     = Conv_out[665];
    assign  image_1_163[15:0]      = Conv_out[664];

    assign  image_1_164[143:128]   = Conv_out[725];
    assign  image_1_164[127:112]   = Conv_out[724];
    assign  image_1_164[111:96]    = Conv_out[723];
    assign  image_1_164[95:80]     = Conv_out[695];
    assign  image_1_164[79:64]     = Conv_out[694];
    assign  image_1_164[63:48]     = Conv_out[693];
    assign  image_1_164[47:32]     = Conv_out[665];
    assign  image_1_164[31:16]     = Conv_out[664];
    assign  image_1_164[15:0]      = Conv_out[663];

    assign  image_1_165[143:128]   = Conv_out[724];
    assign  image_1_165[127:112]   = Conv_out[723];
    assign  image_1_165[111:96]    = Conv_out[722];
    assign  image_1_165[95:80]     = Conv_out[694];
    assign  image_1_165[79:64]     = Conv_out[693];
    assign  image_1_165[63:48]     = Conv_out[692];
    assign  image_1_165[47:32]     = Conv_out[664];
    assign  image_1_165[31:16]     = Conv_out[663];
    assign  image_1_165[15:0]      = Conv_out[662];

    assign  image_1_166[143:128]   = Conv_out[723];
    assign  image_1_166[127:112]   = Conv_out[722];
    assign  image_1_166[111:96]    = Conv_out[721];
    assign  image_1_166[95:80]     = Conv_out[693];
    assign  image_1_166[79:64]     = Conv_out[692];
    assign  image_1_166[63:48]     = Conv_out[691];
    assign  image_1_166[47:32]     = Conv_out[663];
    assign  image_1_166[31:16]     = Conv_out[662];
    assign  image_1_166[15:0]      = Conv_out[661];

    assign  image_1_167[143:128]   = Conv_out[722];
    assign  image_1_167[127:112]   = Conv_out[721];
    assign  image_1_167[111:96]    = Conv_out[720];
    assign  image_1_167[95:80]     = Conv_out[692];
    assign  image_1_167[79:64]     = Conv_out[691];
    assign  image_1_167[63:48]     = Conv_out[690];
    assign  image_1_167[47:32]     = Conv_out[662];
    assign  image_1_167[31:16]     = Conv_out[661];
    assign  image_1_167[15:0]      = Conv_out[660];

    assign  image_1_168[143:128]   = Conv_out[719];
    assign  image_1_168[127:112]   = Conv_out[718];
    assign  image_1_168[111:96]    = Conv_out[717];
    assign  image_1_168[95:80]     = Conv_out[689];
    assign  image_1_168[79:64]     = Conv_out[688];
    assign  image_1_168[63:48]     = Conv_out[687];
    assign  image_1_168[47:32]     = Conv_out[659];
    assign  image_1_168[31:16]     = Conv_out[658];
    assign  image_1_168[15:0]      = Conv_out[657];

    assign  image_1_169[143:128]   = Conv_out[718];
    assign  image_1_169[127:112]   = Conv_out[717];
    assign  image_1_169[111:96]    = Conv_out[716];
    assign  image_1_169[95:80]     = Conv_out[688];
    assign  image_1_169[79:64]     = Conv_out[687];
    assign  image_1_169[63:48]     = Conv_out[686];
    assign  image_1_169[47:32]     = Conv_out[658];
    assign  image_1_169[31:16]     = Conv_out[657];
    assign  image_1_169[15:0]      = Conv_out[656];

    assign  image_1_170[143:128]   = Conv_out[717];
    assign  image_1_170[127:112]   = Conv_out[716];
    assign  image_1_170[111:96]    = Conv_out[715];
    assign  image_1_170[95:80]     = Conv_out[687];
    assign  image_1_170[79:64]     = Conv_out[686];
    assign  image_1_170[63:48]     = Conv_out[685];
    assign  image_1_170[47:32]     = Conv_out[657];
    assign  image_1_170[31:16]     = Conv_out[656];
    assign  image_1_170[15:0]      = Conv_out[655];

    assign  image_1_171[143:128]   = Conv_out[716];
    assign  image_1_171[127:112]   = Conv_out[715];
    assign  image_1_171[111:96]    = Conv_out[714];
    assign  image_1_171[95:80]     = Conv_out[686];
    assign  image_1_171[79:64]     = Conv_out[685];
    assign  image_1_171[63:48]     = Conv_out[684];
    assign  image_1_171[47:32]     = Conv_out[656];
    assign  image_1_171[31:16]     = Conv_out[655];
    assign  image_1_171[15:0]      = Conv_out[654];

    assign  image_1_172[143:128]   = Conv_out[715];
    assign  image_1_172[127:112]   = Conv_out[714];
    assign  image_1_172[111:96]    = Conv_out[713];
    assign  image_1_172[95:80]     = Conv_out[685];
    assign  image_1_172[79:64]     = Conv_out[684];
    assign  image_1_172[63:48]     = Conv_out[683];
    assign  image_1_172[47:32]     = Conv_out[655];
    assign  image_1_172[31:16]     = Conv_out[654];
    assign  image_1_172[15:0]      = Conv_out[653];

    assign  image_1_173[143:128]   = Conv_out[714];
    assign  image_1_173[127:112]   = Conv_out[713];
    assign  image_1_173[111:96]    = Conv_out[712];
    assign  image_1_173[95:80]     = Conv_out[684];
    assign  image_1_173[79:64]     = Conv_out[683];
    assign  image_1_173[63:48]     = Conv_out[682];
    assign  image_1_173[47:32]     = Conv_out[654];
    assign  image_1_173[31:16]     = Conv_out[653];
    assign  image_1_173[15:0]      = Conv_out[652];

    assign  image_1_174[143:128]   = Conv_out[713];
    assign  image_1_174[127:112]   = Conv_out[712];
    assign  image_1_174[111:96]    = Conv_out[711];
    assign  image_1_174[95:80]     = Conv_out[683];
    assign  image_1_174[79:64]     = Conv_out[682];
    assign  image_1_174[63:48]     = Conv_out[681];
    assign  image_1_174[47:32]     = Conv_out[653];
    assign  image_1_174[31:16]     = Conv_out[652];
    assign  image_1_174[15:0]      = Conv_out[651];

    assign  image_1_175[143:128]   = Conv_out[712];
    assign  image_1_175[127:112]   = Conv_out[711];
    assign  image_1_175[111:96]    = Conv_out[710];
    assign  image_1_175[95:80]     = Conv_out[682];
    assign  image_1_175[79:64]     = Conv_out[681];
    assign  image_1_175[63:48]     = Conv_out[680];
    assign  image_1_175[47:32]     = Conv_out[652];
    assign  image_1_175[31:16]     = Conv_out[651];
    assign  image_1_175[15:0]      = Conv_out[650];

    assign  image_1_176[143:128]   = Conv_out[711];
    assign  image_1_176[127:112]   = Conv_out[710];
    assign  image_1_176[111:96]    = Conv_out[709];
    assign  image_1_176[95:80]     = Conv_out[681];
    assign  image_1_176[79:64]     = Conv_out[680];
    assign  image_1_176[63:48]     = Conv_out[679];
    assign  image_1_176[47:32]     = Conv_out[651];
    assign  image_1_176[31:16]     = Conv_out[650];
    assign  image_1_176[15:0]      = Conv_out[649];

    assign  image_1_177[143:128]   = Conv_out[710];
    assign  image_1_177[127:112]   = Conv_out[709];
    assign  image_1_177[111:96]    = Conv_out[708];
    assign  image_1_177[95:80]     = Conv_out[680];
    assign  image_1_177[79:64]     = Conv_out[679];
    assign  image_1_177[63:48]     = Conv_out[678];
    assign  image_1_177[47:32]     = Conv_out[650];
    assign  image_1_177[31:16]     = Conv_out[649];
    assign  image_1_177[15:0]      = Conv_out[648];

    assign  image_1_178[143:128]   = Conv_out[709];
    assign  image_1_178[127:112]   = Conv_out[708];
    assign  image_1_178[111:96]    = Conv_out[707];
    assign  image_1_178[95:80]     = Conv_out[679];
    assign  image_1_178[79:64]     = Conv_out[678];
    assign  image_1_178[63:48]     = Conv_out[677];
    assign  image_1_178[47:32]     = Conv_out[649];
    assign  image_1_178[31:16]     = Conv_out[648];
    assign  image_1_178[15:0]      = Conv_out[647];

    assign  image_1_179[143:128]   = Conv_out[708];
    assign  image_1_179[127:112]   = Conv_out[707];
    assign  image_1_179[111:96]    = Conv_out[706];
    assign  image_1_179[95:80]     = Conv_out[678];
    assign  image_1_179[79:64]     = Conv_out[677];
    assign  image_1_179[63:48]     = Conv_out[676];
    assign  image_1_179[47:32]     = Conv_out[648];
    assign  image_1_179[31:16]     = Conv_out[647];
    assign  image_1_179[15:0]      = Conv_out[646];

    assign  image_1_180[143:128]   = Conv_out[707];
    assign  image_1_180[127:112]   = Conv_out[706];
    assign  image_1_180[111:96]    = Conv_out[705];
    assign  image_1_180[95:80]     = Conv_out[677];
    assign  image_1_180[79:64]     = Conv_out[676];
    assign  image_1_180[63:48]     = Conv_out[675];
    assign  image_1_180[47:32]     = Conv_out[647];
    assign  image_1_180[31:16]     = Conv_out[646];
    assign  image_1_180[15:0]      = Conv_out[645];

    assign  image_1_181[143:128]   = Conv_out[706];
    assign  image_1_181[127:112]   = Conv_out[705];
    assign  image_1_181[111:96]    = Conv_out[704];
    assign  image_1_181[95:80]     = Conv_out[676];
    assign  image_1_181[79:64]     = Conv_out[675];
    assign  image_1_181[63:48]     = Conv_out[674];
    assign  image_1_181[47:32]     = Conv_out[646];
    assign  image_1_181[31:16]     = Conv_out[645];
    assign  image_1_181[15:0]      = Conv_out[644];

    assign  image_1_182[143:128]   = Conv_out[705];
    assign  image_1_182[127:112]   = Conv_out[704];
    assign  image_1_182[111:96]    = Conv_out[703];
    assign  image_1_182[95:80]     = Conv_out[675];
    assign  image_1_182[79:64]     = Conv_out[674];
    assign  image_1_182[63:48]     = Conv_out[673];
    assign  image_1_182[47:32]     = Conv_out[645];
    assign  image_1_182[31:16]     = Conv_out[644];
    assign  image_1_182[15:0]      = Conv_out[643];

    assign  image_1_183[143:128]   = Conv_out[704];
    assign  image_1_183[127:112]   = Conv_out[703];
    assign  image_1_183[111:96]    = Conv_out[702];
    assign  image_1_183[95:80]     = Conv_out[674];
    assign  image_1_183[79:64]     = Conv_out[673];
    assign  image_1_183[63:48]     = Conv_out[672];
    assign  image_1_183[47:32]     = Conv_out[644];
    assign  image_1_183[31:16]     = Conv_out[643];
    assign  image_1_183[15:0]      = Conv_out[642];

    assign  image_1_184[143:128]   = Conv_out[703];
    assign  image_1_184[127:112]   = Conv_out[702];
    assign  image_1_184[111:96]    = Conv_out[701];
    assign  image_1_184[95:80]     = Conv_out[673];
    assign  image_1_184[79:64]     = Conv_out[672];
    assign  image_1_184[63:48]     = Conv_out[671];
    assign  image_1_184[47:32]     = Conv_out[643];
    assign  image_1_184[31:16]     = Conv_out[642];
    assign  image_1_184[15:0]      = Conv_out[641];

    assign  image_1_185[143:128]   = Conv_out[702];
    assign  image_1_185[127:112]   = Conv_out[701];
    assign  image_1_185[111:96]    = Conv_out[700];
    assign  image_1_185[95:80]     = Conv_out[672];
    assign  image_1_185[79:64]     = Conv_out[671];
    assign  image_1_185[63:48]     = Conv_out[670];
    assign  image_1_185[47:32]     = Conv_out[642];
    assign  image_1_185[31:16]     = Conv_out[641];
    assign  image_1_185[15:0]      = Conv_out[640];

    assign  image_1_186[143:128]   = Conv_out[701];
    assign  image_1_186[127:112]   = Conv_out[700];
    assign  image_1_186[111:96]    = Conv_out[699];
    assign  image_1_186[95:80]     = Conv_out[671];
    assign  image_1_186[79:64]     = Conv_out[670];
    assign  image_1_186[63:48]     = Conv_out[669];
    assign  image_1_186[47:32]     = Conv_out[641];
    assign  image_1_186[31:16]     = Conv_out[640];
    assign  image_1_186[15:0]      = Conv_out[639];

    assign  image_1_187[143:128]   = Conv_out[700];
    assign  image_1_187[127:112]   = Conv_out[699];
    assign  image_1_187[111:96]    = Conv_out[698];
    assign  image_1_187[95:80]     = Conv_out[670];
    assign  image_1_187[79:64]     = Conv_out[669];
    assign  image_1_187[63:48]     = Conv_out[668];
    assign  image_1_187[47:32]     = Conv_out[640];
    assign  image_1_187[31:16]     = Conv_out[639];
    assign  image_1_187[15:0]      = Conv_out[638];

    assign  image_1_188[143:128]   = Conv_out[699];
    assign  image_1_188[127:112]   = Conv_out[698];
    assign  image_1_188[111:96]    = Conv_out[697];
    assign  image_1_188[95:80]     = Conv_out[669];
    assign  image_1_188[79:64]     = Conv_out[668];
    assign  image_1_188[63:48]     = Conv_out[667];
    assign  image_1_188[47:32]     = Conv_out[639];
    assign  image_1_188[31:16]     = Conv_out[638];
    assign  image_1_188[15:0]      = Conv_out[637];

    assign  image_1_189[143:128]   = Conv_out[698];
    assign  image_1_189[127:112]   = Conv_out[697];
    assign  image_1_189[111:96]    = Conv_out[696];
    assign  image_1_189[95:80]     = Conv_out[668];
    assign  image_1_189[79:64]     = Conv_out[667];
    assign  image_1_189[63:48]     = Conv_out[666];
    assign  image_1_189[47:32]     = Conv_out[638];
    assign  image_1_189[31:16]     = Conv_out[637];
    assign  image_1_189[15:0]      = Conv_out[636];

    assign  image_1_190[143:128]   = Conv_out[697];
    assign  image_1_190[127:112]   = Conv_out[696];
    assign  image_1_190[111:96]    = Conv_out[695];
    assign  image_1_190[95:80]     = Conv_out[667];
    assign  image_1_190[79:64]     = Conv_out[666];
    assign  image_1_190[63:48]     = Conv_out[665];
    assign  image_1_190[47:32]     = Conv_out[637];
    assign  image_1_190[31:16]     = Conv_out[636];
    assign  image_1_190[15:0]      = Conv_out[635];

    assign  image_1_191[143:128]   = Conv_out[696];
    assign  image_1_191[127:112]   = Conv_out[695];
    assign  image_1_191[111:96]    = Conv_out[694];
    assign  image_1_191[95:80]     = Conv_out[666];
    assign  image_1_191[79:64]     = Conv_out[665];
    assign  image_1_191[63:48]     = Conv_out[664];
    assign  image_1_191[47:32]     = Conv_out[636];
    assign  image_1_191[31:16]     = Conv_out[635];
    assign  image_1_191[15:0]      = Conv_out[634];

    assign  image_1_192[143:128]   = Conv_out[695];
    assign  image_1_192[127:112]   = Conv_out[694];
    assign  image_1_192[111:96]    = Conv_out[693];
    assign  image_1_192[95:80]     = Conv_out[665];
    assign  image_1_192[79:64]     = Conv_out[664];
    assign  image_1_192[63:48]     = Conv_out[663];
    assign  image_1_192[47:32]     = Conv_out[635];
    assign  image_1_192[31:16]     = Conv_out[634];
    assign  image_1_192[15:0]      = Conv_out[633];

    assign  image_1_193[143:128]   = Conv_out[694];
    assign  image_1_193[127:112]   = Conv_out[693];
    assign  image_1_193[111:96]    = Conv_out[692];
    assign  image_1_193[95:80]     = Conv_out[664];
    assign  image_1_193[79:64]     = Conv_out[663];
    assign  image_1_193[63:48]     = Conv_out[662];
    assign  image_1_193[47:32]     = Conv_out[634];
    assign  image_1_193[31:16]     = Conv_out[633];
    assign  image_1_193[15:0]      = Conv_out[632];

    assign  image_1_194[143:128]   = Conv_out[693];
    assign  image_1_194[127:112]   = Conv_out[692];
    assign  image_1_194[111:96]    = Conv_out[691];
    assign  image_1_194[95:80]     = Conv_out[663];
    assign  image_1_194[79:64]     = Conv_out[662];
    assign  image_1_194[63:48]     = Conv_out[661];
    assign  image_1_194[47:32]     = Conv_out[633];
    assign  image_1_194[31:16]     = Conv_out[632];
    assign  image_1_194[15:0]      = Conv_out[631];

    assign  image_1_195[143:128]   = Conv_out[692];
    assign  image_1_195[127:112]   = Conv_out[691];
    assign  image_1_195[111:96]    = Conv_out[690];
    assign  image_1_195[95:80]     = Conv_out[662];
    assign  image_1_195[79:64]     = Conv_out[661];
    assign  image_1_195[63:48]     = Conv_out[660];
    assign  image_1_195[47:32]     = Conv_out[632];
    assign  image_1_195[31:16]     = Conv_out[631];
    assign  image_1_195[15:0]      = Conv_out[630];

    assign  image_1_196[143:128]   = Conv_out[689];
    assign  image_1_196[127:112]   = Conv_out[688];
    assign  image_1_196[111:96]    = Conv_out[687];
    assign  image_1_196[95:80]     = Conv_out[659];
    assign  image_1_196[79:64]     = Conv_out[658];
    assign  image_1_196[63:48]     = Conv_out[657];
    assign  image_1_196[47:32]     = Conv_out[629];
    assign  image_1_196[31:16]     = Conv_out[628];
    assign  image_1_196[15:0]      = Conv_out[627];

    assign  image_1_197[143:128]   = Conv_out[688];
    assign  image_1_197[127:112]   = Conv_out[687];
    assign  image_1_197[111:96]    = Conv_out[686];
    assign  image_1_197[95:80]     = Conv_out[658];
    assign  image_1_197[79:64]     = Conv_out[657];
    assign  image_1_197[63:48]     = Conv_out[656];
    assign  image_1_197[47:32]     = Conv_out[628];
    assign  image_1_197[31:16]     = Conv_out[627];
    assign  image_1_197[15:0]      = Conv_out[626];

    assign  image_1_198[143:128]   = Conv_out[687];
    assign  image_1_198[127:112]   = Conv_out[686];
    assign  image_1_198[111:96]    = Conv_out[685];
    assign  image_1_198[95:80]     = Conv_out[657];
    assign  image_1_198[79:64]     = Conv_out[656];
    assign  image_1_198[63:48]     = Conv_out[655];
    assign  image_1_198[47:32]     = Conv_out[627];
    assign  image_1_198[31:16]     = Conv_out[626];
    assign  image_1_198[15:0]      = Conv_out[625];

    assign  image_1_199[143:128]   = Conv_out[686];
    assign  image_1_199[127:112]   = Conv_out[685];
    assign  image_1_199[111:96]    = Conv_out[684];
    assign  image_1_199[95:80]     = Conv_out[656];
    assign  image_1_199[79:64]     = Conv_out[655];
    assign  image_1_199[63:48]     = Conv_out[654];
    assign  image_1_199[47:32]     = Conv_out[626];
    assign  image_1_199[31:16]     = Conv_out[625];
    assign  image_1_199[15:0]      = Conv_out[624];

    assign  image_1_200[143:128]   = Conv_out[685];
    assign  image_1_200[127:112]   = Conv_out[684];
    assign  image_1_200[111:96]    = Conv_out[683];
    assign  image_1_200[95:80]     = Conv_out[655];
    assign  image_1_200[79:64]     = Conv_out[654];
    assign  image_1_200[63:48]     = Conv_out[653];
    assign  image_1_200[47:32]     = Conv_out[625];
    assign  image_1_200[31:16]     = Conv_out[624];
    assign  image_1_200[15:0]      = Conv_out[623];

    assign  image_1_201[143:128]   = Conv_out[684];
    assign  image_1_201[127:112]   = Conv_out[683];
    assign  image_1_201[111:96]    = Conv_out[682];
    assign  image_1_201[95:80]     = Conv_out[654];
    assign  image_1_201[79:64]     = Conv_out[653];
    assign  image_1_201[63:48]     = Conv_out[652];
    assign  image_1_201[47:32]     = Conv_out[624];
    assign  image_1_201[31:16]     = Conv_out[623];
    assign  image_1_201[15:0]      = Conv_out[622];

    assign  image_1_202[143:128]   = Conv_out[683];
    assign  image_1_202[127:112]   = Conv_out[682];
    assign  image_1_202[111:96]    = Conv_out[681];
    assign  image_1_202[95:80]     = Conv_out[653];
    assign  image_1_202[79:64]     = Conv_out[652];
    assign  image_1_202[63:48]     = Conv_out[651];
    assign  image_1_202[47:32]     = Conv_out[623];
    assign  image_1_202[31:16]     = Conv_out[622];
    assign  image_1_202[15:0]      = Conv_out[621];

    assign  image_1_203[143:128]   = Conv_out[682];
    assign  image_1_203[127:112]   = Conv_out[681];
    assign  image_1_203[111:96]    = Conv_out[680];
    assign  image_1_203[95:80]     = Conv_out[652];
    assign  image_1_203[79:64]     = Conv_out[651];
    assign  image_1_203[63:48]     = Conv_out[650];
    assign  image_1_203[47:32]     = Conv_out[622];
    assign  image_1_203[31:16]     = Conv_out[621];
    assign  image_1_203[15:0]      = Conv_out[620];

    assign  image_1_204[143:128]   = Conv_out[681];
    assign  image_1_204[127:112]   = Conv_out[680];
    assign  image_1_204[111:96]    = Conv_out[679];
    assign  image_1_204[95:80]     = Conv_out[651];
    assign  image_1_204[79:64]     = Conv_out[650];
    assign  image_1_204[63:48]     = Conv_out[649];
    assign  image_1_204[47:32]     = Conv_out[621];
    assign  image_1_204[31:16]     = Conv_out[620];
    assign  image_1_204[15:0]      = Conv_out[619];

    assign  image_1_205[143:128]   = Conv_out[680];
    assign  image_1_205[127:112]   = Conv_out[679];
    assign  image_1_205[111:96]    = Conv_out[678];
    assign  image_1_205[95:80]     = Conv_out[650];
    assign  image_1_205[79:64]     = Conv_out[649];
    assign  image_1_205[63:48]     = Conv_out[648];
    assign  image_1_205[47:32]     = Conv_out[620];
    assign  image_1_205[31:16]     = Conv_out[619];
    assign  image_1_205[15:0]      = Conv_out[618];

    assign  image_1_206[143:128]   = Conv_out[679];
    assign  image_1_206[127:112]   = Conv_out[678];
    assign  image_1_206[111:96]    = Conv_out[677];
    assign  image_1_206[95:80]     = Conv_out[649];
    assign  image_1_206[79:64]     = Conv_out[648];
    assign  image_1_206[63:48]     = Conv_out[647];
    assign  image_1_206[47:32]     = Conv_out[619];
    assign  image_1_206[31:16]     = Conv_out[618];
    assign  image_1_206[15:0]      = Conv_out[617];

    assign  image_1_207[143:128]   = Conv_out[678];
    assign  image_1_207[127:112]   = Conv_out[677];
    assign  image_1_207[111:96]    = Conv_out[676];
    assign  image_1_207[95:80]     = Conv_out[648];
    assign  image_1_207[79:64]     = Conv_out[647];
    assign  image_1_207[63:48]     = Conv_out[646];
    assign  image_1_207[47:32]     = Conv_out[618];
    assign  image_1_207[31:16]     = Conv_out[617];
    assign  image_1_207[15:0]      = Conv_out[616];

    assign  image_1_208[143:128]   = Conv_out[677];
    assign  image_1_208[127:112]   = Conv_out[676];
    assign  image_1_208[111:96]    = Conv_out[675];
    assign  image_1_208[95:80]     = Conv_out[647];
    assign  image_1_208[79:64]     = Conv_out[646];
    assign  image_1_208[63:48]     = Conv_out[645];
    assign  image_1_208[47:32]     = Conv_out[617];
    assign  image_1_208[31:16]     = Conv_out[616];
    assign  image_1_208[15:0]      = Conv_out[615];

    assign  image_1_209[143:128]   = Conv_out[676];
    assign  image_1_209[127:112]   = Conv_out[675];
    assign  image_1_209[111:96]    = Conv_out[674];
    assign  image_1_209[95:80]     = Conv_out[646];
    assign  image_1_209[79:64]     = Conv_out[645];
    assign  image_1_209[63:48]     = Conv_out[644];
    assign  image_1_209[47:32]     = Conv_out[616];
    assign  image_1_209[31:16]     = Conv_out[615];
    assign  image_1_209[15:0]      = Conv_out[614];

    assign  image_1_210[143:128]   = Conv_out[675];
    assign  image_1_210[127:112]   = Conv_out[674];
    assign  image_1_210[111:96]    = Conv_out[673];
    assign  image_1_210[95:80]     = Conv_out[645];
    assign  image_1_210[79:64]     = Conv_out[644];
    assign  image_1_210[63:48]     = Conv_out[643];
    assign  image_1_210[47:32]     = Conv_out[615];
    assign  image_1_210[31:16]     = Conv_out[614];
    assign  image_1_210[15:0]      = Conv_out[613];

    assign  image_1_211[143:128]   = Conv_out[674];
    assign  image_1_211[127:112]   = Conv_out[673];
    assign  image_1_211[111:96]    = Conv_out[672];
    assign  image_1_211[95:80]     = Conv_out[644];
    assign  image_1_211[79:64]     = Conv_out[643];
    assign  image_1_211[63:48]     = Conv_out[642];
    assign  image_1_211[47:32]     = Conv_out[614];
    assign  image_1_211[31:16]     = Conv_out[613];
    assign  image_1_211[15:0]      = Conv_out[612];

    assign  image_1_212[143:128]   = Conv_out[673];
    assign  image_1_212[127:112]   = Conv_out[672];
    assign  image_1_212[111:96]    = Conv_out[671];
    assign  image_1_212[95:80]     = Conv_out[643];
    assign  image_1_212[79:64]     = Conv_out[642];
    assign  image_1_212[63:48]     = Conv_out[641];
    assign  image_1_212[47:32]     = Conv_out[613];
    assign  image_1_212[31:16]     = Conv_out[612];
    assign  image_1_212[15:0]      = Conv_out[611];

    assign  image_1_213[143:128]   = Conv_out[672];
    assign  image_1_213[127:112]   = Conv_out[671];
    assign  image_1_213[111:96]    = Conv_out[670];
    assign  image_1_213[95:80]     = Conv_out[642];
    assign  image_1_213[79:64]     = Conv_out[641];
    assign  image_1_213[63:48]     = Conv_out[640];
    assign  image_1_213[47:32]     = Conv_out[612];
    assign  image_1_213[31:16]     = Conv_out[611];
    assign  image_1_213[15:0]      = Conv_out[610];

    assign  image_1_214[143:128]   = Conv_out[671];
    assign  image_1_214[127:112]   = Conv_out[670];
    assign  image_1_214[111:96]    = Conv_out[669];
    assign  image_1_214[95:80]     = Conv_out[641];
    assign  image_1_214[79:64]     = Conv_out[640];
    assign  image_1_214[63:48]     = Conv_out[639];
    assign  image_1_214[47:32]     = Conv_out[611];
    assign  image_1_214[31:16]     = Conv_out[610];
    assign  image_1_214[15:0]      = Conv_out[609];

    assign  image_1_215[143:128]   = Conv_out[670];
    assign  image_1_215[127:112]   = Conv_out[669];
    assign  image_1_215[111:96]    = Conv_out[668];
    assign  image_1_215[95:80]     = Conv_out[640];
    assign  image_1_215[79:64]     = Conv_out[639];
    assign  image_1_215[63:48]     = Conv_out[638];
    assign  image_1_215[47:32]     = Conv_out[610];
    assign  image_1_215[31:16]     = Conv_out[609];
    assign  image_1_215[15:0]      = Conv_out[608];

    assign  image_1_216[143:128]   = Conv_out[669];
    assign  image_1_216[127:112]   = Conv_out[668];
    assign  image_1_216[111:96]    = Conv_out[667];
    assign  image_1_216[95:80]     = Conv_out[639];
    assign  image_1_216[79:64]     = Conv_out[638];
    assign  image_1_216[63:48]     = Conv_out[637];
    assign  image_1_216[47:32]     = Conv_out[609];
    assign  image_1_216[31:16]     = Conv_out[608];
    assign  image_1_216[15:0]      = Conv_out[607];

    assign  image_1_217[143:128]   = Conv_out[668];
    assign  image_1_217[127:112]   = Conv_out[667];
    assign  image_1_217[111:96]    = Conv_out[666];
    assign  image_1_217[95:80]     = Conv_out[638];
    assign  image_1_217[79:64]     = Conv_out[637];
    assign  image_1_217[63:48]     = Conv_out[636];
    assign  image_1_217[47:32]     = Conv_out[608];
    assign  image_1_217[31:16]     = Conv_out[607];
    assign  image_1_217[15:0]      = Conv_out[606];

    assign  image_1_218[143:128]   = Conv_out[667];
    assign  image_1_218[127:112]   = Conv_out[666];
    assign  image_1_218[111:96]    = Conv_out[665];
    assign  image_1_218[95:80]     = Conv_out[637];
    assign  image_1_218[79:64]     = Conv_out[636];
    assign  image_1_218[63:48]     = Conv_out[635];
    assign  image_1_218[47:32]     = Conv_out[607];
    assign  image_1_218[31:16]     = Conv_out[606];
    assign  image_1_218[15:0]      = Conv_out[605];

    assign  image_1_219[143:128]   = Conv_out[666];
    assign  image_1_219[127:112]   = Conv_out[665];
    assign  image_1_219[111:96]    = Conv_out[664];
    assign  image_1_219[95:80]     = Conv_out[636];
    assign  image_1_219[79:64]     = Conv_out[635];
    assign  image_1_219[63:48]     = Conv_out[634];
    assign  image_1_219[47:32]     = Conv_out[606];
    assign  image_1_219[31:16]     = Conv_out[605];
    assign  image_1_219[15:0]      = Conv_out[604];

    assign  image_1_220[143:128]   = Conv_out[665];
    assign  image_1_220[127:112]   = Conv_out[664];
    assign  image_1_220[111:96]    = Conv_out[663];
    assign  image_1_220[95:80]     = Conv_out[635];
    assign  image_1_220[79:64]     = Conv_out[634];
    assign  image_1_220[63:48]     = Conv_out[633];
    assign  image_1_220[47:32]     = Conv_out[605];
    assign  image_1_220[31:16]     = Conv_out[604];
    assign  image_1_220[15:0]      = Conv_out[603];

    assign  image_1_221[143:128]   = Conv_out[664];
    assign  image_1_221[127:112]   = Conv_out[663];
    assign  image_1_221[111:96]    = Conv_out[662];
    assign  image_1_221[95:80]     = Conv_out[634];
    assign  image_1_221[79:64]     = Conv_out[633];
    assign  image_1_221[63:48]     = Conv_out[632];
    assign  image_1_221[47:32]     = Conv_out[604];
    assign  image_1_221[31:16]     = Conv_out[603];
    assign  image_1_221[15:0]      = Conv_out[602];

    assign  image_1_222[143:128]   = Conv_out[663];
    assign  image_1_222[127:112]   = Conv_out[662];
    assign  image_1_222[111:96]    = Conv_out[661];
    assign  image_1_222[95:80]     = Conv_out[633];
    assign  image_1_222[79:64]     = Conv_out[632];
    assign  image_1_222[63:48]     = Conv_out[631];
    assign  image_1_222[47:32]     = Conv_out[603];
    assign  image_1_222[31:16]     = Conv_out[602];
    assign  image_1_222[15:0]      = Conv_out[601];

    assign  image_1_223[143:128]   = Conv_out[662];
    assign  image_1_223[127:112]   = Conv_out[661];
    assign  image_1_223[111:96]    = Conv_out[660];
    assign  image_1_223[95:80]     = Conv_out[632];
    assign  image_1_223[79:64]     = Conv_out[631];
    assign  image_1_223[63:48]     = Conv_out[630];
    assign  image_1_223[47:32]     = Conv_out[602];
    assign  image_1_223[31:16]     = Conv_out[601];
    assign  image_1_223[15:0]      = Conv_out[600];

    assign  image_1_224[143:128]   = Conv_out[659];
    assign  image_1_224[127:112]   = Conv_out[658];
    assign  image_1_224[111:96]    = Conv_out[657];
    assign  image_1_224[95:80]     = Conv_out[629];
    assign  image_1_224[79:64]     = Conv_out[628];
    assign  image_1_224[63:48]     = Conv_out[627];
    assign  image_1_224[47:32]     = Conv_out[599];
    assign  image_1_224[31:16]     = Conv_out[598];
    assign  image_1_224[15:0]      = Conv_out[597];

    assign  image_1_225[143:128]   = Conv_out[658];
    assign  image_1_225[127:112]   = Conv_out[657];
    assign  image_1_225[111:96]    = Conv_out[656];
    assign  image_1_225[95:80]     = Conv_out[628];
    assign  image_1_225[79:64]     = Conv_out[627];
    assign  image_1_225[63:48]     = Conv_out[626];
    assign  image_1_225[47:32]     = Conv_out[598];
    assign  image_1_225[31:16]     = Conv_out[597];
    assign  image_1_225[15:0]      = Conv_out[596];

    assign  image_1_226[143:128]   = Conv_out[657];
    assign  image_1_226[127:112]   = Conv_out[656];
    assign  image_1_226[111:96]    = Conv_out[655];
    assign  image_1_226[95:80]     = Conv_out[627];
    assign  image_1_226[79:64]     = Conv_out[626];
    assign  image_1_226[63:48]     = Conv_out[625];
    assign  image_1_226[47:32]     = Conv_out[597];
    assign  image_1_226[31:16]     = Conv_out[596];
    assign  image_1_226[15:0]      = Conv_out[595];

    assign  image_1_227[143:128]   = Conv_out[656];
    assign  image_1_227[127:112]   = Conv_out[655];
    assign  image_1_227[111:96]    = Conv_out[654];
    assign  image_1_227[95:80]     = Conv_out[626];
    assign  image_1_227[79:64]     = Conv_out[625];
    assign  image_1_227[63:48]     = Conv_out[624];
    assign  image_1_227[47:32]     = Conv_out[596];
    assign  image_1_227[31:16]     = Conv_out[595];
    assign  image_1_227[15:0]      = Conv_out[594];

    assign  image_1_228[143:128]   = Conv_out[655];
    assign  image_1_228[127:112]   = Conv_out[654];
    assign  image_1_228[111:96]    = Conv_out[653];
    assign  image_1_228[95:80]     = Conv_out[625];
    assign  image_1_228[79:64]     = Conv_out[624];
    assign  image_1_228[63:48]     = Conv_out[623];
    assign  image_1_228[47:32]     = Conv_out[595];
    assign  image_1_228[31:16]     = Conv_out[594];
    assign  image_1_228[15:0]      = Conv_out[593];

    assign  image_1_229[143:128]   = Conv_out[654];
    assign  image_1_229[127:112]   = Conv_out[653];
    assign  image_1_229[111:96]    = Conv_out[652];
    assign  image_1_229[95:80]     = Conv_out[624];
    assign  image_1_229[79:64]     = Conv_out[623];
    assign  image_1_229[63:48]     = Conv_out[622];
    assign  image_1_229[47:32]     = Conv_out[594];
    assign  image_1_229[31:16]     = Conv_out[593];
    assign  image_1_229[15:0]      = Conv_out[592];

    assign  image_1_230[143:128]   = Conv_out[653];
    assign  image_1_230[127:112]   = Conv_out[652];
    assign  image_1_230[111:96]    = Conv_out[651];
    assign  image_1_230[95:80]     = Conv_out[623];
    assign  image_1_230[79:64]     = Conv_out[622];
    assign  image_1_230[63:48]     = Conv_out[621];
    assign  image_1_230[47:32]     = Conv_out[593];
    assign  image_1_230[31:16]     = Conv_out[592];
    assign  image_1_230[15:0]      = Conv_out[591];

    assign  image_1_231[143:128]   = Conv_out[652];
    assign  image_1_231[127:112]   = Conv_out[651];
    assign  image_1_231[111:96]    = Conv_out[650];
    assign  image_1_231[95:80]     = Conv_out[622];
    assign  image_1_231[79:64]     = Conv_out[621];
    assign  image_1_231[63:48]     = Conv_out[620];
    assign  image_1_231[47:32]     = Conv_out[592];
    assign  image_1_231[31:16]     = Conv_out[591];
    assign  image_1_231[15:0]      = Conv_out[590];

    assign  image_1_232[143:128]   = Conv_out[651];
    assign  image_1_232[127:112]   = Conv_out[650];
    assign  image_1_232[111:96]    = Conv_out[649];
    assign  image_1_232[95:80]     = Conv_out[621];
    assign  image_1_232[79:64]     = Conv_out[620];
    assign  image_1_232[63:48]     = Conv_out[619];
    assign  image_1_232[47:32]     = Conv_out[591];
    assign  image_1_232[31:16]     = Conv_out[590];
    assign  image_1_232[15:0]      = Conv_out[589];

    assign  image_1_233[143:128]   = Conv_out[650];
    assign  image_1_233[127:112]   = Conv_out[649];
    assign  image_1_233[111:96]    = Conv_out[648];
    assign  image_1_233[95:80]     = Conv_out[620];
    assign  image_1_233[79:64]     = Conv_out[619];
    assign  image_1_233[63:48]     = Conv_out[618];
    assign  image_1_233[47:32]     = Conv_out[590];
    assign  image_1_233[31:16]     = Conv_out[589];
    assign  image_1_233[15:0]      = Conv_out[588];

    assign  image_1_234[143:128]   = Conv_out[649];
    assign  image_1_234[127:112]   = Conv_out[648];
    assign  image_1_234[111:96]    = Conv_out[647];
    assign  image_1_234[95:80]     = Conv_out[619];
    assign  image_1_234[79:64]     = Conv_out[618];
    assign  image_1_234[63:48]     = Conv_out[617];
    assign  image_1_234[47:32]     = Conv_out[589];
    assign  image_1_234[31:16]     = Conv_out[588];
    assign  image_1_234[15:0]      = Conv_out[587];

    assign  image_1_235[143:128]   = Conv_out[648];
    assign  image_1_235[127:112]   = Conv_out[647];
    assign  image_1_235[111:96]    = Conv_out[646];
    assign  image_1_235[95:80]     = Conv_out[618];
    assign  image_1_235[79:64]     = Conv_out[617];
    assign  image_1_235[63:48]     = Conv_out[616];
    assign  image_1_235[47:32]     = Conv_out[588];
    assign  image_1_235[31:16]     = Conv_out[587];
    assign  image_1_235[15:0]      = Conv_out[586];

    assign  image_1_236[143:128]   = Conv_out[647];
    assign  image_1_236[127:112]   = Conv_out[646];
    assign  image_1_236[111:96]    = Conv_out[645];
    assign  image_1_236[95:80]     = Conv_out[617];
    assign  image_1_236[79:64]     = Conv_out[616];
    assign  image_1_236[63:48]     = Conv_out[615];
    assign  image_1_236[47:32]     = Conv_out[587];
    assign  image_1_236[31:16]     = Conv_out[586];
    assign  image_1_236[15:0]      = Conv_out[585];

    assign  image_1_237[143:128]   = Conv_out[646];
    assign  image_1_237[127:112]   = Conv_out[645];
    assign  image_1_237[111:96]    = Conv_out[644];
    assign  image_1_237[95:80]     = Conv_out[616];
    assign  image_1_237[79:64]     = Conv_out[615];
    assign  image_1_237[63:48]     = Conv_out[614];
    assign  image_1_237[47:32]     = Conv_out[586];
    assign  image_1_237[31:16]     = Conv_out[585];
    assign  image_1_237[15:0]      = Conv_out[584];

    assign  image_1_238[143:128]   = Conv_out[645];
    assign  image_1_238[127:112]   = Conv_out[644];
    assign  image_1_238[111:96]    = Conv_out[643];
    assign  image_1_238[95:80]     = Conv_out[615];
    assign  image_1_238[79:64]     = Conv_out[614];
    assign  image_1_238[63:48]     = Conv_out[613];
    assign  image_1_238[47:32]     = Conv_out[585];
    assign  image_1_238[31:16]     = Conv_out[584];
    assign  image_1_238[15:0]      = Conv_out[583];

    assign  image_1_239[143:128]   = Conv_out[644];
    assign  image_1_239[127:112]   = Conv_out[643];
    assign  image_1_239[111:96]    = Conv_out[642];
    assign  image_1_239[95:80]     = Conv_out[614];
    assign  image_1_239[79:64]     = Conv_out[613];
    assign  image_1_239[63:48]     = Conv_out[612];
    assign  image_1_239[47:32]     = Conv_out[584];
    assign  image_1_239[31:16]     = Conv_out[583];
    assign  image_1_239[15:0]      = Conv_out[582];

    assign  image_1_240[143:128]   = Conv_out[643];
    assign  image_1_240[127:112]   = Conv_out[642];
    assign  image_1_240[111:96]    = Conv_out[641];
    assign  image_1_240[95:80]     = Conv_out[613];
    assign  image_1_240[79:64]     = Conv_out[612];
    assign  image_1_240[63:48]     = Conv_out[611];
    assign  image_1_240[47:32]     = Conv_out[583];
    assign  image_1_240[31:16]     = Conv_out[582];
    assign  image_1_240[15:0]      = Conv_out[581];

    assign  image_1_241[143:128]   = Conv_out[642];
    assign  image_1_241[127:112]   = Conv_out[641];
    assign  image_1_241[111:96]    = Conv_out[640];
    assign  image_1_241[95:80]     = Conv_out[612];
    assign  image_1_241[79:64]     = Conv_out[611];
    assign  image_1_241[63:48]     = Conv_out[610];
    assign  image_1_241[47:32]     = Conv_out[582];
    assign  image_1_241[31:16]     = Conv_out[581];
    assign  image_1_241[15:0]      = Conv_out[580];

    assign  image_1_242[143:128]   = Conv_out[641];
    assign  image_1_242[127:112]   = Conv_out[640];
    assign  image_1_242[111:96]    = Conv_out[639];
    assign  image_1_242[95:80]     = Conv_out[611];
    assign  image_1_242[79:64]     = Conv_out[610];
    assign  image_1_242[63:48]     = Conv_out[609];
    assign  image_1_242[47:32]     = Conv_out[581];
    assign  image_1_242[31:16]     = Conv_out[580];
    assign  image_1_242[15:0]      = Conv_out[579];

    assign  image_1_243[143:128]   = Conv_out[640];
    assign  image_1_243[127:112]   = Conv_out[639];
    assign  image_1_243[111:96]    = Conv_out[638];
    assign  image_1_243[95:80]     = Conv_out[610];
    assign  image_1_243[79:64]     = Conv_out[609];
    assign  image_1_243[63:48]     = Conv_out[608];
    assign  image_1_243[47:32]     = Conv_out[580];
    assign  image_1_243[31:16]     = Conv_out[579];
    assign  image_1_243[15:0]      = Conv_out[578];

    assign  image_1_244[143:128]   = Conv_out[639];
    assign  image_1_244[127:112]   = Conv_out[638];
    assign  image_1_244[111:96]    = Conv_out[637];
    assign  image_1_244[95:80]     = Conv_out[609];
    assign  image_1_244[79:64]     = Conv_out[608];
    assign  image_1_244[63:48]     = Conv_out[607];
    assign  image_1_244[47:32]     = Conv_out[579];
    assign  image_1_244[31:16]     = Conv_out[578];
    assign  image_1_244[15:0]      = Conv_out[577];

    assign  image_1_245[143:128]   = Conv_out[638];
    assign  image_1_245[127:112]   = Conv_out[637];
    assign  image_1_245[111:96]    = Conv_out[636];
    assign  image_1_245[95:80]     = Conv_out[608];
    assign  image_1_245[79:64]     = Conv_out[607];
    assign  image_1_245[63:48]     = Conv_out[606];
    assign  image_1_245[47:32]     = Conv_out[578];
    assign  image_1_245[31:16]     = Conv_out[577];
    assign  image_1_245[15:0]      = Conv_out[576];

    assign  image_1_246[143:128]   = Conv_out[637];
    assign  image_1_246[127:112]   = Conv_out[636];
    assign  image_1_246[111:96]    = Conv_out[635];
    assign  image_1_246[95:80]     = Conv_out[607];
    assign  image_1_246[79:64]     = Conv_out[606];
    assign  image_1_246[63:48]     = Conv_out[605];
    assign  image_1_246[47:32]     = Conv_out[577];
    assign  image_1_246[31:16]     = Conv_out[576];
    assign  image_1_246[15:0]      = Conv_out[575];

    assign  image_1_247[143:128]   = Conv_out[636];
    assign  image_1_247[127:112]   = Conv_out[635];
    assign  image_1_247[111:96]    = Conv_out[634];
    assign  image_1_247[95:80]     = Conv_out[606];
    assign  image_1_247[79:64]     = Conv_out[605];
    assign  image_1_247[63:48]     = Conv_out[604];
    assign  image_1_247[47:32]     = Conv_out[576];
    assign  image_1_247[31:16]     = Conv_out[575];
    assign  image_1_247[15:0]      = Conv_out[574];

    assign  image_1_248[143:128]   = Conv_out[635];
    assign  image_1_248[127:112]   = Conv_out[634];
    assign  image_1_248[111:96]    = Conv_out[633];
    assign  image_1_248[95:80]     = Conv_out[605];
    assign  image_1_248[79:64]     = Conv_out[604];
    assign  image_1_248[63:48]     = Conv_out[603];
    assign  image_1_248[47:32]     = Conv_out[575];
    assign  image_1_248[31:16]     = Conv_out[574];
    assign  image_1_248[15:0]      = Conv_out[573];

    assign  image_1_249[143:128]   = Conv_out[634];
    assign  image_1_249[127:112]   = Conv_out[633];
    assign  image_1_249[111:96]    = Conv_out[632];
    assign  image_1_249[95:80]     = Conv_out[604];
    assign  image_1_249[79:64]     = Conv_out[603];
    assign  image_1_249[63:48]     = Conv_out[602];
    assign  image_1_249[47:32]     = Conv_out[574];
    assign  image_1_249[31:16]     = Conv_out[573];
    assign  image_1_249[15:0]      = Conv_out[572];

    assign  image_1_250[143:128]   = Conv_out[633];
    assign  image_1_250[127:112]   = Conv_out[632];
    assign  image_1_250[111:96]    = Conv_out[631];
    assign  image_1_250[95:80]     = Conv_out[603];
    assign  image_1_250[79:64]     = Conv_out[602];
    assign  image_1_250[63:48]     = Conv_out[601];
    assign  image_1_250[47:32]     = Conv_out[573];
    assign  image_1_250[31:16]     = Conv_out[572];
    assign  image_1_250[15:0]      = Conv_out[571];

    assign  image_1_251[143:128]   = Conv_out[632];
    assign  image_1_251[127:112]   = Conv_out[631];
    assign  image_1_251[111:96]    = Conv_out[630];
    assign  image_1_251[95:80]     = Conv_out[602];
    assign  image_1_251[79:64]     = Conv_out[601];
    assign  image_1_251[63:48]     = Conv_out[600];
    assign  image_1_251[47:32]     = Conv_out[572];
    assign  image_1_251[31:16]     = Conv_out[571];
    assign  image_1_251[15:0]      = Conv_out[570];

    assign  image_1_252[143:128]   = Conv_out[629];
    assign  image_1_252[127:112]   = Conv_out[628];
    assign  image_1_252[111:96]    = Conv_out[627];
    assign  image_1_252[95:80]     = Conv_out[599];
    assign  image_1_252[79:64]     = Conv_out[598];
    assign  image_1_252[63:48]     = Conv_out[597];
    assign  image_1_252[47:32]     = Conv_out[569];
    assign  image_1_252[31:16]     = Conv_out[568];
    assign  image_1_252[15:0]      = Conv_out[567];

    assign  image_1_253[143:128]   = Conv_out[628];
    assign  image_1_253[127:112]   = Conv_out[627];
    assign  image_1_253[111:96]    = Conv_out[626];
    assign  image_1_253[95:80]     = Conv_out[598];
    assign  image_1_253[79:64]     = Conv_out[597];
    assign  image_1_253[63:48]     = Conv_out[596];
    assign  image_1_253[47:32]     = Conv_out[568];
    assign  image_1_253[31:16]     = Conv_out[567];
    assign  image_1_253[15:0]      = Conv_out[566];

    assign  image_1_254[143:128]   = Conv_out[627];
    assign  image_1_254[127:112]   = Conv_out[626];
    assign  image_1_254[111:96]    = Conv_out[625];
    assign  image_1_254[95:80]     = Conv_out[597];
    assign  image_1_254[79:64]     = Conv_out[596];
    assign  image_1_254[63:48]     = Conv_out[595];
    assign  image_1_254[47:32]     = Conv_out[567];
    assign  image_1_254[31:16]     = Conv_out[566];
    assign  image_1_254[15:0]      = Conv_out[565];

    assign  image_1_255[143:128]   = Conv_out[626];
    assign  image_1_255[127:112]   = Conv_out[625];
    assign  image_1_255[111:96]    = Conv_out[624];
    assign  image_1_255[95:80]     = Conv_out[596];
    assign  image_1_255[79:64]     = Conv_out[595];
    assign  image_1_255[63:48]     = Conv_out[594];
    assign  image_1_255[47:32]     = Conv_out[566];
    assign  image_1_255[31:16]     = Conv_out[565];
    assign  image_1_255[15:0]      = Conv_out[564];

    assign  image_1_256[143:128]   = Conv_out[625];
    assign  image_1_256[127:112]   = Conv_out[624];
    assign  image_1_256[111:96]    = Conv_out[623];
    assign  image_1_256[95:80]     = Conv_out[595];
    assign  image_1_256[79:64]     = Conv_out[594];
    assign  image_1_256[63:48]     = Conv_out[593];
    assign  image_1_256[47:32]     = Conv_out[565];
    assign  image_1_256[31:16]     = Conv_out[564];
    assign  image_1_256[15:0]      = Conv_out[563];

    assign  image_1_257[143:128]   = Conv_out[624];
    assign  image_1_257[127:112]   = Conv_out[623];
    assign  image_1_257[111:96]    = Conv_out[622];
    assign  image_1_257[95:80]     = Conv_out[594];
    assign  image_1_257[79:64]     = Conv_out[593];
    assign  image_1_257[63:48]     = Conv_out[592];
    assign  image_1_257[47:32]     = Conv_out[564];
    assign  image_1_257[31:16]     = Conv_out[563];
    assign  image_1_257[15:0]      = Conv_out[562];

    assign  image_1_258[143:128]   = Conv_out[623];
    assign  image_1_258[127:112]   = Conv_out[622];
    assign  image_1_258[111:96]    = Conv_out[621];
    assign  image_1_258[95:80]     = Conv_out[593];
    assign  image_1_258[79:64]     = Conv_out[592];
    assign  image_1_258[63:48]     = Conv_out[591];
    assign  image_1_258[47:32]     = Conv_out[563];
    assign  image_1_258[31:16]     = Conv_out[562];
    assign  image_1_258[15:0]      = Conv_out[561];

    assign  image_1_259[143:128]   = Conv_out[622];
    assign  image_1_259[127:112]   = Conv_out[621];
    assign  image_1_259[111:96]    = Conv_out[620];
    assign  image_1_259[95:80]     = Conv_out[592];
    assign  image_1_259[79:64]     = Conv_out[591];
    assign  image_1_259[63:48]     = Conv_out[590];
    assign  image_1_259[47:32]     = Conv_out[562];
    assign  image_1_259[31:16]     = Conv_out[561];
    assign  image_1_259[15:0]      = Conv_out[560];

    assign  image_1_260[143:128]   = Conv_out[621];
    assign  image_1_260[127:112]   = Conv_out[620];
    assign  image_1_260[111:96]    = Conv_out[619];
    assign  image_1_260[95:80]     = Conv_out[591];
    assign  image_1_260[79:64]     = Conv_out[590];
    assign  image_1_260[63:48]     = Conv_out[589];
    assign  image_1_260[47:32]     = Conv_out[561];
    assign  image_1_260[31:16]     = Conv_out[560];
    assign  image_1_260[15:0]      = Conv_out[559];

    assign  image_1_261[143:128]   = Conv_out[620];
    assign  image_1_261[127:112]   = Conv_out[619];
    assign  image_1_261[111:96]    = Conv_out[618];
    assign  image_1_261[95:80]     = Conv_out[590];
    assign  image_1_261[79:64]     = Conv_out[589];
    assign  image_1_261[63:48]     = Conv_out[588];
    assign  image_1_261[47:32]     = Conv_out[560];
    assign  image_1_261[31:16]     = Conv_out[559];
    assign  image_1_261[15:0]      = Conv_out[558];

    assign  image_1_262[143:128]   = Conv_out[619];
    assign  image_1_262[127:112]   = Conv_out[618];
    assign  image_1_262[111:96]    = Conv_out[617];
    assign  image_1_262[95:80]     = Conv_out[589];
    assign  image_1_262[79:64]     = Conv_out[588];
    assign  image_1_262[63:48]     = Conv_out[587];
    assign  image_1_262[47:32]     = Conv_out[559];
    assign  image_1_262[31:16]     = Conv_out[558];
    assign  image_1_262[15:0]      = Conv_out[557];

    assign  image_1_263[143:128]   = Conv_out[618];
    assign  image_1_263[127:112]   = Conv_out[617];
    assign  image_1_263[111:96]    = Conv_out[616];
    assign  image_1_263[95:80]     = Conv_out[588];
    assign  image_1_263[79:64]     = Conv_out[587];
    assign  image_1_263[63:48]     = Conv_out[586];
    assign  image_1_263[47:32]     = Conv_out[558];
    assign  image_1_263[31:16]     = Conv_out[557];
    assign  image_1_263[15:0]      = Conv_out[556];

    assign  image_1_264[143:128]   = Conv_out[617];
    assign  image_1_264[127:112]   = Conv_out[616];
    assign  image_1_264[111:96]    = Conv_out[615];
    assign  image_1_264[95:80]     = Conv_out[587];
    assign  image_1_264[79:64]     = Conv_out[586];
    assign  image_1_264[63:48]     = Conv_out[585];
    assign  image_1_264[47:32]     = Conv_out[557];
    assign  image_1_264[31:16]     = Conv_out[556];
    assign  image_1_264[15:0]      = Conv_out[555];

    assign  image_1_265[143:128]   = Conv_out[616];
    assign  image_1_265[127:112]   = Conv_out[615];
    assign  image_1_265[111:96]    = Conv_out[614];
    assign  image_1_265[95:80]     = Conv_out[586];
    assign  image_1_265[79:64]     = Conv_out[585];
    assign  image_1_265[63:48]     = Conv_out[584];
    assign  image_1_265[47:32]     = Conv_out[556];
    assign  image_1_265[31:16]     = Conv_out[555];
    assign  image_1_265[15:0]      = Conv_out[554];

    assign  image_1_266[143:128]   = Conv_out[615];
    assign  image_1_266[127:112]   = Conv_out[614];
    assign  image_1_266[111:96]    = Conv_out[613];
    assign  image_1_266[95:80]     = Conv_out[585];
    assign  image_1_266[79:64]     = Conv_out[584];
    assign  image_1_266[63:48]     = Conv_out[583];
    assign  image_1_266[47:32]     = Conv_out[555];
    assign  image_1_266[31:16]     = Conv_out[554];
    assign  image_1_266[15:0]      = Conv_out[553];

    assign  image_1_267[143:128]   = Conv_out[614];
    assign  image_1_267[127:112]   = Conv_out[613];
    assign  image_1_267[111:96]    = Conv_out[612];
    assign  image_1_267[95:80]     = Conv_out[584];
    assign  image_1_267[79:64]     = Conv_out[583];
    assign  image_1_267[63:48]     = Conv_out[582];
    assign  image_1_267[47:32]     = Conv_out[554];
    assign  image_1_267[31:16]     = Conv_out[553];
    assign  image_1_267[15:0]      = Conv_out[552];

    assign  image_1_268[143:128]   = Conv_out[613];
    assign  image_1_268[127:112]   = Conv_out[612];
    assign  image_1_268[111:96]    = Conv_out[611];
    assign  image_1_268[95:80]     = Conv_out[583];
    assign  image_1_268[79:64]     = Conv_out[582];
    assign  image_1_268[63:48]     = Conv_out[581];
    assign  image_1_268[47:32]     = Conv_out[553];
    assign  image_1_268[31:16]     = Conv_out[552];
    assign  image_1_268[15:0]      = Conv_out[551];

    assign  image_1_269[143:128]   = Conv_out[612];
    assign  image_1_269[127:112]   = Conv_out[611];
    assign  image_1_269[111:96]    = Conv_out[610];
    assign  image_1_269[95:80]     = Conv_out[582];
    assign  image_1_269[79:64]     = Conv_out[581];
    assign  image_1_269[63:48]     = Conv_out[580];
    assign  image_1_269[47:32]     = Conv_out[552];
    assign  image_1_269[31:16]     = Conv_out[551];
    assign  image_1_269[15:0]      = Conv_out[550];

    assign  image_1_270[143:128]   = Conv_out[611];
    assign  image_1_270[127:112]   = Conv_out[610];
    assign  image_1_270[111:96]    = Conv_out[609];
    assign  image_1_270[95:80]     = Conv_out[581];
    assign  image_1_270[79:64]     = Conv_out[580];
    assign  image_1_270[63:48]     = Conv_out[579];
    assign  image_1_270[47:32]     = Conv_out[551];
    assign  image_1_270[31:16]     = Conv_out[550];
    assign  image_1_270[15:0]      = Conv_out[549];

    assign  image_1_271[143:128]   = Conv_out[610];
    assign  image_1_271[127:112]   = Conv_out[609];
    assign  image_1_271[111:96]    = Conv_out[608];
    assign  image_1_271[95:80]     = Conv_out[580];
    assign  image_1_271[79:64]     = Conv_out[579];
    assign  image_1_271[63:48]     = Conv_out[578];
    assign  image_1_271[47:32]     = Conv_out[550];
    assign  image_1_271[31:16]     = Conv_out[549];
    assign  image_1_271[15:0]      = Conv_out[548];

    assign  image_1_272[143:128]   = Conv_out[609];
    assign  image_1_272[127:112]   = Conv_out[608];
    assign  image_1_272[111:96]    = Conv_out[607];
    assign  image_1_272[95:80]     = Conv_out[579];
    assign  image_1_272[79:64]     = Conv_out[578];
    assign  image_1_272[63:48]     = Conv_out[577];
    assign  image_1_272[47:32]     = Conv_out[549];
    assign  image_1_272[31:16]     = Conv_out[548];
    assign  image_1_272[15:0]      = Conv_out[547];

    assign  image_1_273[143:128]   = Conv_out[608];
    assign  image_1_273[127:112]   = Conv_out[607];
    assign  image_1_273[111:96]    = Conv_out[606];
    assign  image_1_273[95:80]     = Conv_out[578];
    assign  image_1_273[79:64]     = Conv_out[577];
    assign  image_1_273[63:48]     = Conv_out[576];
    assign  image_1_273[47:32]     = Conv_out[548];
    assign  image_1_273[31:16]     = Conv_out[547];
    assign  image_1_273[15:0]      = Conv_out[546];

    assign  image_1_274[143:128]   = Conv_out[607];
    assign  image_1_274[127:112]   = Conv_out[606];
    assign  image_1_274[111:96]    = Conv_out[605];
    assign  image_1_274[95:80]     = Conv_out[577];
    assign  image_1_274[79:64]     = Conv_out[576];
    assign  image_1_274[63:48]     = Conv_out[575];
    assign  image_1_274[47:32]     = Conv_out[547];
    assign  image_1_274[31:16]     = Conv_out[546];
    assign  image_1_274[15:0]      = Conv_out[545];

    assign  image_1_275[143:128]   = Conv_out[606];
    assign  image_1_275[127:112]   = Conv_out[605];
    assign  image_1_275[111:96]    = Conv_out[604];
    assign  image_1_275[95:80]     = Conv_out[576];
    assign  image_1_275[79:64]     = Conv_out[575];
    assign  image_1_275[63:48]     = Conv_out[574];
    assign  image_1_275[47:32]     = Conv_out[546];
    assign  image_1_275[31:16]     = Conv_out[545];
    assign  image_1_275[15:0]      = Conv_out[544];

    assign  image_1_276[143:128]   = Conv_out[605];
    assign  image_1_276[127:112]   = Conv_out[604];
    assign  image_1_276[111:96]    = Conv_out[603];
    assign  image_1_276[95:80]     = Conv_out[575];
    assign  image_1_276[79:64]     = Conv_out[574];
    assign  image_1_276[63:48]     = Conv_out[573];
    assign  image_1_276[47:32]     = Conv_out[545];
    assign  image_1_276[31:16]     = Conv_out[544];
    assign  image_1_276[15:0]      = Conv_out[543];

    assign  image_1_277[143:128]   = Conv_out[604];
    assign  image_1_277[127:112]   = Conv_out[603];
    assign  image_1_277[111:96]    = Conv_out[602];
    assign  image_1_277[95:80]     = Conv_out[574];
    assign  image_1_277[79:64]     = Conv_out[573];
    assign  image_1_277[63:48]     = Conv_out[572];
    assign  image_1_277[47:32]     = Conv_out[544];
    assign  image_1_277[31:16]     = Conv_out[543];
    assign  image_1_277[15:0]      = Conv_out[542];

    assign  image_1_278[143:128]   = Conv_out[603];
    assign  image_1_278[127:112]   = Conv_out[602];
    assign  image_1_278[111:96]    = Conv_out[601];
    assign  image_1_278[95:80]     = Conv_out[573];
    assign  image_1_278[79:64]     = Conv_out[572];
    assign  image_1_278[63:48]     = Conv_out[571];
    assign  image_1_278[47:32]     = Conv_out[543];
    assign  image_1_278[31:16]     = Conv_out[542];
    assign  image_1_278[15:0]      = Conv_out[541];

    assign  image_1_279[143:128]   = Conv_out[602];
    assign  image_1_279[127:112]   = Conv_out[601];
    assign  image_1_279[111:96]    = Conv_out[600];
    assign  image_1_279[95:80]     = Conv_out[572];
    assign  image_1_279[79:64]     = Conv_out[571];
    assign  image_1_279[63:48]     = Conv_out[570];
    assign  image_1_279[47:32]     = Conv_out[542];
    assign  image_1_279[31:16]     = Conv_out[541];
    assign  image_1_279[15:0]      = Conv_out[540];

    assign  image_1_280[143:128]   = Conv_out[599];
    assign  image_1_280[127:112]   = Conv_out[598];
    assign  image_1_280[111:96]    = Conv_out[597];
    assign  image_1_280[95:80]     = Conv_out[569];
    assign  image_1_280[79:64]     = Conv_out[568];
    assign  image_1_280[63:48]     = Conv_out[567];
    assign  image_1_280[47:32]     = Conv_out[539];
    assign  image_1_280[31:16]     = Conv_out[538];
    assign  image_1_280[15:0]      = Conv_out[537];

    assign  image_1_281[143:128]   = Conv_out[598];
    assign  image_1_281[127:112]   = Conv_out[597];
    assign  image_1_281[111:96]    = Conv_out[596];
    assign  image_1_281[95:80]     = Conv_out[568];
    assign  image_1_281[79:64]     = Conv_out[567];
    assign  image_1_281[63:48]     = Conv_out[566];
    assign  image_1_281[47:32]     = Conv_out[538];
    assign  image_1_281[31:16]     = Conv_out[537];
    assign  image_1_281[15:0]      = Conv_out[536];

    assign  image_1_282[143:128]   = Conv_out[597];
    assign  image_1_282[127:112]   = Conv_out[596];
    assign  image_1_282[111:96]    = Conv_out[595];
    assign  image_1_282[95:80]     = Conv_out[567];
    assign  image_1_282[79:64]     = Conv_out[566];
    assign  image_1_282[63:48]     = Conv_out[565];
    assign  image_1_282[47:32]     = Conv_out[537];
    assign  image_1_282[31:16]     = Conv_out[536];
    assign  image_1_282[15:0]      = Conv_out[535];

    assign  image_1_283[143:128]   = Conv_out[596];
    assign  image_1_283[127:112]   = Conv_out[595];
    assign  image_1_283[111:96]    = Conv_out[594];
    assign  image_1_283[95:80]     = Conv_out[566];
    assign  image_1_283[79:64]     = Conv_out[565];
    assign  image_1_283[63:48]     = Conv_out[564];
    assign  image_1_283[47:32]     = Conv_out[536];
    assign  image_1_283[31:16]     = Conv_out[535];
    assign  image_1_283[15:0]      = Conv_out[534];

    assign  image_1_284[143:128]   = Conv_out[595];
    assign  image_1_284[127:112]   = Conv_out[594];
    assign  image_1_284[111:96]    = Conv_out[593];
    assign  image_1_284[95:80]     = Conv_out[565];
    assign  image_1_284[79:64]     = Conv_out[564];
    assign  image_1_284[63:48]     = Conv_out[563];
    assign  image_1_284[47:32]     = Conv_out[535];
    assign  image_1_284[31:16]     = Conv_out[534];
    assign  image_1_284[15:0]      = Conv_out[533];

    assign  image_1_285[143:128]   = Conv_out[594];
    assign  image_1_285[127:112]   = Conv_out[593];
    assign  image_1_285[111:96]    = Conv_out[592];
    assign  image_1_285[95:80]     = Conv_out[564];
    assign  image_1_285[79:64]     = Conv_out[563];
    assign  image_1_285[63:48]     = Conv_out[562];
    assign  image_1_285[47:32]     = Conv_out[534];
    assign  image_1_285[31:16]     = Conv_out[533];
    assign  image_1_285[15:0]      = Conv_out[532];

    assign  image_1_286[143:128]   = Conv_out[593];
    assign  image_1_286[127:112]   = Conv_out[592];
    assign  image_1_286[111:96]    = Conv_out[591];
    assign  image_1_286[95:80]     = Conv_out[563];
    assign  image_1_286[79:64]     = Conv_out[562];
    assign  image_1_286[63:48]     = Conv_out[561];
    assign  image_1_286[47:32]     = Conv_out[533];
    assign  image_1_286[31:16]     = Conv_out[532];
    assign  image_1_286[15:0]      = Conv_out[531];

    assign  image_1_287[143:128]   = Conv_out[592];
    assign  image_1_287[127:112]   = Conv_out[591];
    assign  image_1_287[111:96]    = Conv_out[590];
    assign  image_1_287[95:80]     = Conv_out[562];
    assign  image_1_287[79:64]     = Conv_out[561];
    assign  image_1_287[63:48]     = Conv_out[560];
    assign  image_1_287[47:32]     = Conv_out[532];
    assign  image_1_287[31:16]     = Conv_out[531];
    assign  image_1_287[15:0]      = Conv_out[530];

    assign  image_1_288[143:128]   = Conv_out[591];
    assign  image_1_288[127:112]   = Conv_out[590];
    assign  image_1_288[111:96]    = Conv_out[589];
    assign  image_1_288[95:80]     = Conv_out[561];
    assign  image_1_288[79:64]     = Conv_out[560];
    assign  image_1_288[63:48]     = Conv_out[559];
    assign  image_1_288[47:32]     = Conv_out[531];
    assign  image_1_288[31:16]     = Conv_out[530];
    assign  image_1_288[15:0]      = Conv_out[529];

    assign  image_1_289[143:128]   = Conv_out[590];
    assign  image_1_289[127:112]   = Conv_out[589];
    assign  image_1_289[111:96]    = Conv_out[588];
    assign  image_1_289[95:80]     = Conv_out[560];
    assign  image_1_289[79:64]     = Conv_out[559];
    assign  image_1_289[63:48]     = Conv_out[558];
    assign  image_1_289[47:32]     = Conv_out[530];
    assign  image_1_289[31:16]     = Conv_out[529];
    assign  image_1_289[15:0]      = Conv_out[528];

    assign  image_1_290[143:128]   = Conv_out[589];
    assign  image_1_290[127:112]   = Conv_out[588];
    assign  image_1_290[111:96]    = Conv_out[587];
    assign  image_1_290[95:80]     = Conv_out[559];
    assign  image_1_290[79:64]     = Conv_out[558];
    assign  image_1_290[63:48]     = Conv_out[557];
    assign  image_1_290[47:32]     = Conv_out[529];
    assign  image_1_290[31:16]     = Conv_out[528];
    assign  image_1_290[15:0]      = Conv_out[527];

    assign  image_1_291[143:128]   = Conv_out[588];
    assign  image_1_291[127:112]   = Conv_out[587];
    assign  image_1_291[111:96]    = Conv_out[586];
    assign  image_1_291[95:80]     = Conv_out[558];
    assign  image_1_291[79:64]     = Conv_out[557];
    assign  image_1_291[63:48]     = Conv_out[556];
    assign  image_1_291[47:32]     = Conv_out[528];
    assign  image_1_291[31:16]     = Conv_out[527];
    assign  image_1_291[15:0]      = Conv_out[526];

    assign  image_1_292[143:128]   = Conv_out[587];
    assign  image_1_292[127:112]   = Conv_out[586];
    assign  image_1_292[111:96]    = Conv_out[585];
    assign  image_1_292[95:80]     = Conv_out[557];
    assign  image_1_292[79:64]     = Conv_out[556];
    assign  image_1_292[63:48]     = Conv_out[555];
    assign  image_1_292[47:32]     = Conv_out[527];
    assign  image_1_292[31:16]     = Conv_out[526];
    assign  image_1_292[15:0]      = Conv_out[525];

    assign  image_1_293[143:128]   = Conv_out[586];
    assign  image_1_293[127:112]   = Conv_out[585];
    assign  image_1_293[111:96]    = Conv_out[584];
    assign  image_1_293[95:80]     = Conv_out[556];
    assign  image_1_293[79:64]     = Conv_out[555];
    assign  image_1_293[63:48]     = Conv_out[554];
    assign  image_1_293[47:32]     = Conv_out[526];
    assign  image_1_293[31:16]     = Conv_out[525];
    assign  image_1_293[15:0]      = Conv_out[524];

    assign  image_1_294[143:128]   = Conv_out[585];
    assign  image_1_294[127:112]   = Conv_out[584];
    assign  image_1_294[111:96]    = Conv_out[583];
    assign  image_1_294[95:80]     = Conv_out[555];
    assign  image_1_294[79:64]     = Conv_out[554];
    assign  image_1_294[63:48]     = Conv_out[553];
    assign  image_1_294[47:32]     = Conv_out[525];
    assign  image_1_294[31:16]     = Conv_out[524];
    assign  image_1_294[15:0]      = Conv_out[523];

    assign  image_1_295[143:128]   = Conv_out[584];
    assign  image_1_295[127:112]   = Conv_out[583];
    assign  image_1_295[111:96]    = Conv_out[582];
    assign  image_1_295[95:80]     = Conv_out[554];
    assign  image_1_295[79:64]     = Conv_out[553];
    assign  image_1_295[63:48]     = Conv_out[552];
    assign  image_1_295[47:32]     = Conv_out[524];
    assign  image_1_295[31:16]     = Conv_out[523];
    assign  image_1_295[15:0]      = Conv_out[522];

    assign  image_1_296[143:128]   = Conv_out[583];
    assign  image_1_296[127:112]   = Conv_out[582];
    assign  image_1_296[111:96]    = Conv_out[581];
    assign  image_1_296[95:80]     = Conv_out[553];
    assign  image_1_296[79:64]     = Conv_out[552];
    assign  image_1_296[63:48]     = Conv_out[551];
    assign  image_1_296[47:32]     = Conv_out[523];
    assign  image_1_296[31:16]     = Conv_out[522];
    assign  image_1_296[15:0]      = Conv_out[521];

    assign  image_1_297[143:128]   = Conv_out[582];
    assign  image_1_297[127:112]   = Conv_out[581];
    assign  image_1_297[111:96]    = Conv_out[580];
    assign  image_1_297[95:80]     = Conv_out[552];
    assign  image_1_297[79:64]     = Conv_out[551];
    assign  image_1_297[63:48]     = Conv_out[550];
    assign  image_1_297[47:32]     = Conv_out[522];
    assign  image_1_297[31:16]     = Conv_out[521];
    assign  image_1_297[15:0]      = Conv_out[520];

    assign  image_1_298[143:128]   = Conv_out[581];
    assign  image_1_298[127:112]   = Conv_out[580];
    assign  image_1_298[111:96]    = Conv_out[579];
    assign  image_1_298[95:80]     = Conv_out[551];
    assign  image_1_298[79:64]     = Conv_out[550];
    assign  image_1_298[63:48]     = Conv_out[549];
    assign  image_1_298[47:32]     = Conv_out[521];
    assign  image_1_298[31:16]     = Conv_out[520];
    assign  image_1_298[15:0]      = Conv_out[519];

    assign  image_1_299[143:128]   = Conv_out[580];
    assign  image_1_299[127:112]   = Conv_out[579];
    assign  image_1_299[111:96]    = Conv_out[578];
    assign  image_1_299[95:80]     = Conv_out[550];
    assign  image_1_299[79:64]     = Conv_out[549];
    assign  image_1_299[63:48]     = Conv_out[548];
    assign  image_1_299[47:32]     = Conv_out[520];
    assign  image_1_299[31:16]     = Conv_out[519];
    assign  image_1_299[15:0]      = Conv_out[518];

    assign  image_1_300[143:128]   = Conv_out[579];
    assign  image_1_300[127:112]   = Conv_out[578];
    assign  image_1_300[111:96]    = Conv_out[577];
    assign  image_1_300[95:80]     = Conv_out[549];
    assign  image_1_300[79:64]     = Conv_out[548];
    assign  image_1_300[63:48]     = Conv_out[547];
    assign  image_1_300[47:32]     = Conv_out[519];
    assign  image_1_300[31:16]     = Conv_out[518];
    assign  image_1_300[15:0]      = Conv_out[517];

    assign  image_1_301[143:128]   = Conv_out[578];
    assign  image_1_301[127:112]   = Conv_out[577];
    assign  image_1_301[111:96]    = Conv_out[576];
    assign  image_1_301[95:80]     = Conv_out[548];
    assign  image_1_301[79:64]     = Conv_out[547];
    assign  image_1_301[63:48]     = Conv_out[546];
    assign  image_1_301[47:32]     = Conv_out[518];
    assign  image_1_301[31:16]     = Conv_out[517];
    assign  image_1_301[15:0]      = Conv_out[516];

    assign  image_1_302[143:128]   = Conv_out[577];
    assign  image_1_302[127:112]   = Conv_out[576];
    assign  image_1_302[111:96]    = Conv_out[575];
    assign  image_1_302[95:80]     = Conv_out[547];
    assign  image_1_302[79:64]     = Conv_out[546];
    assign  image_1_302[63:48]     = Conv_out[545];
    assign  image_1_302[47:32]     = Conv_out[517];
    assign  image_1_302[31:16]     = Conv_out[516];
    assign  image_1_302[15:0]      = Conv_out[515];

    assign  image_1_303[143:128]   = Conv_out[576];
    assign  image_1_303[127:112]   = Conv_out[575];
    assign  image_1_303[111:96]    = Conv_out[574];
    assign  image_1_303[95:80]     = Conv_out[546];
    assign  image_1_303[79:64]     = Conv_out[545];
    assign  image_1_303[63:48]     = Conv_out[544];
    assign  image_1_303[47:32]     = Conv_out[516];
    assign  image_1_303[31:16]     = Conv_out[515];
    assign  image_1_303[15:0]      = Conv_out[514];

    assign  image_1_304[143:128]   = Conv_out[575];
    assign  image_1_304[127:112]   = Conv_out[574];
    assign  image_1_304[111:96]    = Conv_out[573];
    assign  image_1_304[95:80]     = Conv_out[545];
    assign  image_1_304[79:64]     = Conv_out[544];
    assign  image_1_304[63:48]     = Conv_out[543];
    assign  image_1_304[47:32]     = Conv_out[515];
    assign  image_1_304[31:16]     = Conv_out[514];
    assign  image_1_304[15:0]      = Conv_out[513];

    assign  image_1_305[143:128]   = Conv_out[574];
    assign  image_1_305[127:112]   = Conv_out[573];
    assign  image_1_305[111:96]    = Conv_out[572];
    assign  image_1_305[95:80]     = Conv_out[544];
    assign  image_1_305[79:64]     = Conv_out[543];
    assign  image_1_305[63:48]     = Conv_out[542];
    assign  image_1_305[47:32]     = Conv_out[514];
    assign  image_1_305[31:16]     = Conv_out[513];
    assign  image_1_305[15:0]      = Conv_out[512];

    assign  image_1_306[143:128]   = Conv_out[573];
    assign  image_1_306[127:112]   = Conv_out[572];
    assign  image_1_306[111:96]    = Conv_out[571];
    assign  image_1_306[95:80]     = Conv_out[543];
    assign  image_1_306[79:64]     = Conv_out[542];
    assign  image_1_306[63:48]     = Conv_out[541];
    assign  image_1_306[47:32]     = Conv_out[513];
    assign  image_1_306[31:16]     = Conv_out[512];
    assign  image_1_306[15:0]      = Conv_out[511];

    assign  image_1_307[143:128]   = Conv_out[572];
    assign  image_1_307[127:112]   = Conv_out[571];
    assign  image_1_307[111:96]    = Conv_out[570];
    assign  image_1_307[95:80]     = Conv_out[542];
    assign  image_1_307[79:64]     = Conv_out[541];
    assign  image_1_307[63:48]     = Conv_out[540];
    assign  image_1_307[47:32]     = Conv_out[512];
    assign  image_1_307[31:16]     = Conv_out[511];
    assign  image_1_307[15:0]      = Conv_out[510];

    assign  image_1_308[143:128]   = Conv_out[569];
    assign  image_1_308[127:112]   = Conv_out[568];
    assign  image_1_308[111:96]    = Conv_out[567];
    assign  image_1_308[95:80]     = Conv_out[539];
    assign  image_1_308[79:64]     = Conv_out[538];
    assign  image_1_308[63:48]     = Conv_out[537];
    assign  image_1_308[47:32]     = Conv_out[509];
    assign  image_1_308[31:16]     = Conv_out[508];
    assign  image_1_308[15:0]      = Conv_out[507];

    assign  image_1_309[143:128]   = Conv_out[568];
    assign  image_1_309[127:112]   = Conv_out[567];
    assign  image_1_309[111:96]    = Conv_out[566];
    assign  image_1_309[95:80]     = Conv_out[538];
    assign  image_1_309[79:64]     = Conv_out[537];
    assign  image_1_309[63:48]     = Conv_out[536];
    assign  image_1_309[47:32]     = Conv_out[508];
    assign  image_1_309[31:16]     = Conv_out[507];
    assign  image_1_309[15:0]      = Conv_out[506];

    assign  image_1_310[143:128]   = Conv_out[567];
    assign  image_1_310[127:112]   = Conv_out[566];
    assign  image_1_310[111:96]    = Conv_out[565];
    assign  image_1_310[95:80]     = Conv_out[537];
    assign  image_1_310[79:64]     = Conv_out[536];
    assign  image_1_310[63:48]     = Conv_out[535];
    assign  image_1_310[47:32]     = Conv_out[507];
    assign  image_1_310[31:16]     = Conv_out[506];
    assign  image_1_310[15:0]      = Conv_out[505];

    assign  image_1_311[143:128]   = Conv_out[566];
    assign  image_1_311[127:112]   = Conv_out[565];
    assign  image_1_311[111:96]    = Conv_out[564];
    assign  image_1_311[95:80]     = Conv_out[536];
    assign  image_1_311[79:64]     = Conv_out[535];
    assign  image_1_311[63:48]     = Conv_out[534];
    assign  image_1_311[47:32]     = Conv_out[506];
    assign  image_1_311[31:16]     = Conv_out[505];
    assign  image_1_311[15:0]      = Conv_out[504];

    assign  image_1_312[143:128]   = Conv_out[565];
    assign  image_1_312[127:112]   = Conv_out[564];
    assign  image_1_312[111:96]    = Conv_out[563];
    assign  image_1_312[95:80]     = Conv_out[535];
    assign  image_1_312[79:64]     = Conv_out[534];
    assign  image_1_312[63:48]     = Conv_out[533];
    assign  image_1_312[47:32]     = Conv_out[505];
    assign  image_1_312[31:16]     = Conv_out[504];
    assign  image_1_312[15:0]      = Conv_out[503];

    assign  image_1_313[143:128]   = Conv_out[564];
    assign  image_1_313[127:112]   = Conv_out[563];
    assign  image_1_313[111:96]    = Conv_out[562];
    assign  image_1_313[95:80]     = Conv_out[534];
    assign  image_1_313[79:64]     = Conv_out[533];
    assign  image_1_313[63:48]     = Conv_out[532];
    assign  image_1_313[47:32]     = Conv_out[504];
    assign  image_1_313[31:16]     = Conv_out[503];
    assign  image_1_313[15:0]      = Conv_out[502];

    assign  image_1_314[143:128]   = Conv_out[563];
    assign  image_1_314[127:112]   = Conv_out[562];
    assign  image_1_314[111:96]    = Conv_out[561];
    assign  image_1_314[95:80]     = Conv_out[533];
    assign  image_1_314[79:64]     = Conv_out[532];
    assign  image_1_314[63:48]     = Conv_out[531];
    assign  image_1_314[47:32]     = Conv_out[503];
    assign  image_1_314[31:16]     = Conv_out[502];
    assign  image_1_314[15:0]      = Conv_out[501];

    assign  image_1_315[143:128]   = Conv_out[562];
    assign  image_1_315[127:112]   = Conv_out[561];
    assign  image_1_315[111:96]    = Conv_out[560];
    assign  image_1_315[95:80]     = Conv_out[532];
    assign  image_1_315[79:64]     = Conv_out[531];
    assign  image_1_315[63:48]     = Conv_out[530];
    assign  image_1_315[47:32]     = Conv_out[502];
    assign  image_1_315[31:16]     = Conv_out[501];
    assign  image_1_315[15:0]      = Conv_out[500];

    assign  image_1_316[143:128]   = Conv_out[561];
    assign  image_1_316[127:112]   = Conv_out[560];
    assign  image_1_316[111:96]    = Conv_out[559];
    assign  image_1_316[95:80]     = Conv_out[531];
    assign  image_1_316[79:64]     = Conv_out[530];
    assign  image_1_316[63:48]     = Conv_out[529];
    assign  image_1_316[47:32]     = Conv_out[501];
    assign  image_1_316[31:16]     = Conv_out[500];
    assign  image_1_316[15:0]      = Conv_out[499];

    assign  image_1_317[143:128]   = Conv_out[560];
    assign  image_1_317[127:112]   = Conv_out[559];
    assign  image_1_317[111:96]    = Conv_out[558];
    assign  image_1_317[95:80]     = Conv_out[530];
    assign  image_1_317[79:64]     = Conv_out[529];
    assign  image_1_317[63:48]     = Conv_out[528];
    assign  image_1_317[47:32]     = Conv_out[500];
    assign  image_1_317[31:16]     = Conv_out[499];
    assign  image_1_317[15:0]      = Conv_out[498];

    assign  image_1_318[143:128]   = Conv_out[559];
    assign  image_1_318[127:112]   = Conv_out[558];
    assign  image_1_318[111:96]    = Conv_out[557];
    assign  image_1_318[95:80]     = Conv_out[529];
    assign  image_1_318[79:64]     = Conv_out[528];
    assign  image_1_318[63:48]     = Conv_out[527];
    assign  image_1_318[47:32]     = Conv_out[499];
    assign  image_1_318[31:16]     = Conv_out[498];
    assign  image_1_318[15:0]      = Conv_out[497];

    assign  image_1_319[143:128]   = Conv_out[558];
    assign  image_1_319[127:112]   = Conv_out[557];
    assign  image_1_319[111:96]    = Conv_out[556];
    assign  image_1_319[95:80]     = Conv_out[528];
    assign  image_1_319[79:64]     = Conv_out[527];
    assign  image_1_319[63:48]     = Conv_out[526];
    assign  image_1_319[47:32]     = Conv_out[498];
    assign  image_1_319[31:16]     = Conv_out[497];
    assign  image_1_319[15:0]      = Conv_out[496];

    assign  image_1_320[143:128]   = Conv_out[557];
    assign  image_1_320[127:112]   = Conv_out[556];
    assign  image_1_320[111:96]    = Conv_out[555];
    assign  image_1_320[95:80]     = Conv_out[527];
    assign  image_1_320[79:64]     = Conv_out[526];
    assign  image_1_320[63:48]     = Conv_out[525];
    assign  image_1_320[47:32]     = Conv_out[497];
    assign  image_1_320[31:16]     = Conv_out[496];
    assign  image_1_320[15:0]      = Conv_out[495];

    assign  image_1_321[143:128]   = Conv_out[556];
    assign  image_1_321[127:112]   = Conv_out[555];
    assign  image_1_321[111:96]    = Conv_out[554];
    assign  image_1_321[95:80]     = Conv_out[526];
    assign  image_1_321[79:64]     = Conv_out[525];
    assign  image_1_321[63:48]     = Conv_out[524];
    assign  image_1_321[47:32]     = Conv_out[496];
    assign  image_1_321[31:16]     = Conv_out[495];
    assign  image_1_321[15:0]      = Conv_out[494];

    assign  image_1_322[143:128]   = Conv_out[555];
    assign  image_1_322[127:112]   = Conv_out[554];
    assign  image_1_322[111:96]    = Conv_out[553];
    assign  image_1_322[95:80]     = Conv_out[525];
    assign  image_1_322[79:64]     = Conv_out[524];
    assign  image_1_322[63:48]     = Conv_out[523];
    assign  image_1_322[47:32]     = Conv_out[495];
    assign  image_1_322[31:16]     = Conv_out[494];
    assign  image_1_322[15:0]      = Conv_out[493];

    assign  image_1_323[143:128]   = Conv_out[554];
    assign  image_1_323[127:112]   = Conv_out[553];
    assign  image_1_323[111:96]    = Conv_out[552];
    assign  image_1_323[95:80]     = Conv_out[524];
    assign  image_1_323[79:64]     = Conv_out[523];
    assign  image_1_323[63:48]     = Conv_out[522];
    assign  image_1_323[47:32]     = Conv_out[494];
    assign  image_1_323[31:16]     = Conv_out[493];
    assign  image_1_323[15:0]      = Conv_out[492];

    assign  image_1_324[143:128]   = Conv_out[553];
    assign  image_1_324[127:112]   = Conv_out[552];
    assign  image_1_324[111:96]    = Conv_out[551];
    assign  image_1_324[95:80]     = Conv_out[523];
    assign  image_1_324[79:64]     = Conv_out[522];
    assign  image_1_324[63:48]     = Conv_out[521];
    assign  image_1_324[47:32]     = Conv_out[493];
    assign  image_1_324[31:16]     = Conv_out[492];
    assign  image_1_324[15:0]      = Conv_out[491];

    assign  image_1_325[143:128]   = Conv_out[552];
    assign  image_1_325[127:112]   = Conv_out[551];
    assign  image_1_325[111:96]    = Conv_out[550];
    assign  image_1_325[95:80]     = Conv_out[522];
    assign  image_1_325[79:64]     = Conv_out[521];
    assign  image_1_325[63:48]     = Conv_out[520];
    assign  image_1_325[47:32]     = Conv_out[492];
    assign  image_1_325[31:16]     = Conv_out[491];
    assign  image_1_325[15:0]      = Conv_out[490];

    assign  image_1_326[143:128]   = Conv_out[551];
    assign  image_1_326[127:112]   = Conv_out[550];
    assign  image_1_326[111:96]    = Conv_out[549];
    assign  image_1_326[95:80]     = Conv_out[521];
    assign  image_1_326[79:64]     = Conv_out[520];
    assign  image_1_326[63:48]     = Conv_out[519];
    assign  image_1_326[47:32]     = Conv_out[491];
    assign  image_1_326[31:16]     = Conv_out[490];
    assign  image_1_326[15:0]      = Conv_out[489];

    assign  image_1_327[143:128]   = Conv_out[550];
    assign  image_1_327[127:112]   = Conv_out[549];
    assign  image_1_327[111:96]    = Conv_out[548];
    assign  image_1_327[95:80]     = Conv_out[520];
    assign  image_1_327[79:64]     = Conv_out[519];
    assign  image_1_327[63:48]     = Conv_out[518];
    assign  image_1_327[47:32]     = Conv_out[490];
    assign  image_1_327[31:16]     = Conv_out[489];
    assign  image_1_327[15:0]      = Conv_out[488];

    assign  image_1_328[143:128]   = Conv_out[549];
    assign  image_1_328[127:112]   = Conv_out[548];
    assign  image_1_328[111:96]    = Conv_out[547];
    assign  image_1_328[95:80]     = Conv_out[519];
    assign  image_1_328[79:64]     = Conv_out[518];
    assign  image_1_328[63:48]     = Conv_out[517];
    assign  image_1_328[47:32]     = Conv_out[489];
    assign  image_1_328[31:16]     = Conv_out[488];
    assign  image_1_328[15:0]      = Conv_out[487];

    assign  image_1_329[143:128]   = Conv_out[548];
    assign  image_1_329[127:112]   = Conv_out[547];
    assign  image_1_329[111:96]    = Conv_out[546];
    assign  image_1_329[95:80]     = Conv_out[518];
    assign  image_1_329[79:64]     = Conv_out[517];
    assign  image_1_329[63:48]     = Conv_out[516];
    assign  image_1_329[47:32]     = Conv_out[488];
    assign  image_1_329[31:16]     = Conv_out[487];
    assign  image_1_329[15:0]      = Conv_out[486];

    assign  image_1_330[143:128]   = Conv_out[547];
    assign  image_1_330[127:112]   = Conv_out[546];
    assign  image_1_330[111:96]    = Conv_out[545];
    assign  image_1_330[95:80]     = Conv_out[517];
    assign  image_1_330[79:64]     = Conv_out[516];
    assign  image_1_330[63:48]     = Conv_out[515];
    assign  image_1_330[47:32]     = Conv_out[487];
    assign  image_1_330[31:16]     = Conv_out[486];
    assign  image_1_330[15:0]      = Conv_out[485];

    assign  image_1_331[143:128]   = Conv_out[546];
    assign  image_1_331[127:112]   = Conv_out[545];
    assign  image_1_331[111:96]    = Conv_out[544];
    assign  image_1_331[95:80]     = Conv_out[516];
    assign  image_1_331[79:64]     = Conv_out[515];
    assign  image_1_331[63:48]     = Conv_out[514];
    assign  image_1_331[47:32]     = Conv_out[486];
    assign  image_1_331[31:16]     = Conv_out[485];
    assign  image_1_331[15:0]      = Conv_out[484];

    assign  image_1_332[143:128]   = Conv_out[545];
    assign  image_1_332[127:112]   = Conv_out[544];
    assign  image_1_332[111:96]    = Conv_out[543];
    assign  image_1_332[95:80]     = Conv_out[515];
    assign  image_1_332[79:64]     = Conv_out[514];
    assign  image_1_332[63:48]     = Conv_out[513];
    assign  image_1_332[47:32]     = Conv_out[485];
    assign  image_1_332[31:16]     = Conv_out[484];
    assign  image_1_332[15:0]      = Conv_out[483];

    assign  image_1_333[143:128]   = Conv_out[544];
    assign  image_1_333[127:112]   = Conv_out[543];
    assign  image_1_333[111:96]    = Conv_out[542];
    assign  image_1_333[95:80]     = Conv_out[514];
    assign  image_1_333[79:64]     = Conv_out[513];
    assign  image_1_333[63:48]     = Conv_out[512];
    assign  image_1_333[47:32]     = Conv_out[484];
    assign  image_1_333[31:16]     = Conv_out[483];
    assign  image_1_333[15:0]      = Conv_out[482];

    assign  image_1_334[143:128]   = Conv_out[543];
    assign  image_1_334[127:112]   = Conv_out[542];
    assign  image_1_334[111:96]    = Conv_out[541];
    assign  image_1_334[95:80]     = Conv_out[513];
    assign  image_1_334[79:64]     = Conv_out[512];
    assign  image_1_334[63:48]     = Conv_out[511];
    assign  image_1_334[47:32]     = Conv_out[483];
    assign  image_1_334[31:16]     = Conv_out[482];
    assign  image_1_334[15:0]      = Conv_out[481];

    assign  image_1_335[143:128]   = Conv_out[542];
    assign  image_1_335[127:112]   = Conv_out[541];
    assign  image_1_335[111:96]    = Conv_out[540];
    assign  image_1_335[95:80]     = Conv_out[512];
    assign  image_1_335[79:64]     = Conv_out[511];
    assign  image_1_335[63:48]     = Conv_out[510];
    assign  image_1_335[47:32]     = Conv_out[482];
    assign  image_1_335[31:16]     = Conv_out[481];
    assign  image_1_335[15:0]      = Conv_out[480];

    assign  image_1_336[143:128]   = Conv_out[539];
    assign  image_1_336[127:112]   = Conv_out[538];
    assign  image_1_336[111:96]    = Conv_out[537];
    assign  image_1_336[95:80]     = Conv_out[509];
    assign  image_1_336[79:64]     = Conv_out[508];
    assign  image_1_336[63:48]     = Conv_out[507];
    assign  image_1_336[47:32]     = Conv_out[479];
    assign  image_1_336[31:16]     = Conv_out[478];
    assign  image_1_336[15:0]      = Conv_out[477];

    assign  image_1_337[143:128]   = Conv_out[538];
    assign  image_1_337[127:112]   = Conv_out[537];
    assign  image_1_337[111:96]    = Conv_out[536];
    assign  image_1_337[95:80]     = Conv_out[508];
    assign  image_1_337[79:64]     = Conv_out[507];
    assign  image_1_337[63:48]     = Conv_out[506];
    assign  image_1_337[47:32]     = Conv_out[478];
    assign  image_1_337[31:16]     = Conv_out[477];
    assign  image_1_337[15:0]      = Conv_out[476];

    assign  image_1_338[143:128]   = Conv_out[537];
    assign  image_1_338[127:112]   = Conv_out[536];
    assign  image_1_338[111:96]    = Conv_out[535];
    assign  image_1_338[95:80]     = Conv_out[507];
    assign  image_1_338[79:64]     = Conv_out[506];
    assign  image_1_338[63:48]     = Conv_out[505];
    assign  image_1_338[47:32]     = Conv_out[477];
    assign  image_1_338[31:16]     = Conv_out[476];
    assign  image_1_338[15:0]      = Conv_out[475];

    assign  image_1_339[143:128]   = Conv_out[536];
    assign  image_1_339[127:112]   = Conv_out[535];
    assign  image_1_339[111:96]    = Conv_out[534];
    assign  image_1_339[95:80]     = Conv_out[506];
    assign  image_1_339[79:64]     = Conv_out[505];
    assign  image_1_339[63:48]     = Conv_out[504];
    assign  image_1_339[47:32]     = Conv_out[476];
    assign  image_1_339[31:16]     = Conv_out[475];
    assign  image_1_339[15:0]      = Conv_out[474];

    assign  image_1_340[143:128]   = Conv_out[535];
    assign  image_1_340[127:112]   = Conv_out[534];
    assign  image_1_340[111:96]    = Conv_out[533];
    assign  image_1_340[95:80]     = Conv_out[505];
    assign  image_1_340[79:64]     = Conv_out[504];
    assign  image_1_340[63:48]     = Conv_out[503];
    assign  image_1_340[47:32]     = Conv_out[475];
    assign  image_1_340[31:16]     = Conv_out[474];
    assign  image_1_340[15:0]      = Conv_out[473];

    assign  image_1_341[143:128]   = Conv_out[534];
    assign  image_1_341[127:112]   = Conv_out[533];
    assign  image_1_341[111:96]    = Conv_out[532];
    assign  image_1_341[95:80]     = Conv_out[504];
    assign  image_1_341[79:64]     = Conv_out[503];
    assign  image_1_341[63:48]     = Conv_out[502];
    assign  image_1_341[47:32]     = Conv_out[474];
    assign  image_1_341[31:16]     = Conv_out[473];
    assign  image_1_341[15:0]      = Conv_out[472];

    assign  image_1_342[143:128]   = Conv_out[533];
    assign  image_1_342[127:112]   = Conv_out[532];
    assign  image_1_342[111:96]    = Conv_out[531];
    assign  image_1_342[95:80]     = Conv_out[503];
    assign  image_1_342[79:64]     = Conv_out[502];
    assign  image_1_342[63:48]     = Conv_out[501];
    assign  image_1_342[47:32]     = Conv_out[473];
    assign  image_1_342[31:16]     = Conv_out[472];
    assign  image_1_342[15:0]      = Conv_out[471];

    assign  image_1_343[143:128]   = Conv_out[532];
    assign  image_1_343[127:112]   = Conv_out[531];
    assign  image_1_343[111:96]    = Conv_out[530];
    assign  image_1_343[95:80]     = Conv_out[502];
    assign  image_1_343[79:64]     = Conv_out[501];
    assign  image_1_343[63:48]     = Conv_out[500];
    assign  image_1_343[47:32]     = Conv_out[472];
    assign  image_1_343[31:16]     = Conv_out[471];
    assign  image_1_343[15:0]      = Conv_out[470];

    assign  image_1_344[143:128]   = Conv_out[531];
    assign  image_1_344[127:112]   = Conv_out[530];
    assign  image_1_344[111:96]    = Conv_out[529];
    assign  image_1_344[95:80]     = Conv_out[501];
    assign  image_1_344[79:64]     = Conv_out[500];
    assign  image_1_344[63:48]     = Conv_out[499];
    assign  image_1_344[47:32]     = Conv_out[471];
    assign  image_1_344[31:16]     = Conv_out[470];
    assign  image_1_344[15:0]      = Conv_out[469];

    assign  image_1_345[143:128]   = Conv_out[530];
    assign  image_1_345[127:112]   = Conv_out[529];
    assign  image_1_345[111:96]    = Conv_out[528];
    assign  image_1_345[95:80]     = Conv_out[500];
    assign  image_1_345[79:64]     = Conv_out[499];
    assign  image_1_345[63:48]     = Conv_out[498];
    assign  image_1_345[47:32]     = Conv_out[470];
    assign  image_1_345[31:16]     = Conv_out[469];
    assign  image_1_345[15:0]      = Conv_out[468];

    assign  image_1_346[143:128]   = Conv_out[529];
    assign  image_1_346[127:112]   = Conv_out[528];
    assign  image_1_346[111:96]    = Conv_out[527];
    assign  image_1_346[95:80]     = Conv_out[499];
    assign  image_1_346[79:64]     = Conv_out[498];
    assign  image_1_346[63:48]     = Conv_out[497];
    assign  image_1_346[47:32]     = Conv_out[469];
    assign  image_1_346[31:16]     = Conv_out[468];
    assign  image_1_346[15:0]      = Conv_out[467];

    assign  image_1_347[143:128]   = Conv_out[528];
    assign  image_1_347[127:112]   = Conv_out[527];
    assign  image_1_347[111:96]    = Conv_out[526];
    assign  image_1_347[95:80]     = Conv_out[498];
    assign  image_1_347[79:64]     = Conv_out[497];
    assign  image_1_347[63:48]     = Conv_out[496];
    assign  image_1_347[47:32]     = Conv_out[468];
    assign  image_1_347[31:16]     = Conv_out[467];
    assign  image_1_347[15:0]      = Conv_out[466];

    assign  image_1_348[143:128]   = Conv_out[527];
    assign  image_1_348[127:112]   = Conv_out[526];
    assign  image_1_348[111:96]    = Conv_out[525];
    assign  image_1_348[95:80]     = Conv_out[497];
    assign  image_1_348[79:64]     = Conv_out[496];
    assign  image_1_348[63:48]     = Conv_out[495];
    assign  image_1_348[47:32]     = Conv_out[467];
    assign  image_1_348[31:16]     = Conv_out[466];
    assign  image_1_348[15:0]      = Conv_out[465];

    assign  image_1_349[143:128]   = Conv_out[526];
    assign  image_1_349[127:112]   = Conv_out[525];
    assign  image_1_349[111:96]    = Conv_out[524];
    assign  image_1_349[95:80]     = Conv_out[496];
    assign  image_1_349[79:64]     = Conv_out[495];
    assign  image_1_349[63:48]     = Conv_out[494];
    assign  image_1_349[47:32]     = Conv_out[466];
    assign  image_1_349[31:16]     = Conv_out[465];
    assign  image_1_349[15:0]      = Conv_out[464];

    assign  image_1_350[143:128]   = Conv_out[525];
    assign  image_1_350[127:112]   = Conv_out[524];
    assign  image_1_350[111:96]    = Conv_out[523];
    assign  image_1_350[95:80]     = Conv_out[495];
    assign  image_1_350[79:64]     = Conv_out[494];
    assign  image_1_350[63:48]     = Conv_out[493];
    assign  image_1_350[47:32]     = Conv_out[465];
    assign  image_1_350[31:16]     = Conv_out[464];
    assign  image_1_350[15:0]      = Conv_out[463];

    assign  image_1_351[143:128]   = Conv_out[524];
    assign  image_1_351[127:112]   = Conv_out[523];
    assign  image_1_351[111:96]    = Conv_out[522];
    assign  image_1_351[95:80]     = Conv_out[494];
    assign  image_1_351[79:64]     = Conv_out[493];
    assign  image_1_351[63:48]     = Conv_out[492];
    assign  image_1_351[47:32]     = Conv_out[464];
    assign  image_1_351[31:16]     = Conv_out[463];
    assign  image_1_351[15:0]      = Conv_out[462];

    assign  image_1_352[143:128]   = Conv_out[523];
    assign  image_1_352[127:112]   = Conv_out[522];
    assign  image_1_352[111:96]    = Conv_out[521];
    assign  image_1_352[95:80]     = Conv_out[493];
    assign  image_1_352[79:64]     = Conv_out[492];
    assign  image_1_352[63:48]     = Conv_out[491];
    assign  image_1_352[47:32]     = Conv_out[463];
    assign  image_1_352[31:16]     = Conv_out[462];
    assign  image_1_352[15:0]      = Conv_out[461];

    assign  image_1_353[143:128]   = Conv_out[522];
    assign  image_1_353[127:112]   = Conv_out[521];
    assign  image_1_353[111:96]    = Conv_out[520];
    assign  image_1_353[95:80]     = Conv_out[492];
    assign  image_1_353[79:64]     = Conv_out[491];
    assign  image_1_353[63:48]     = Conv_out[490];
    assign  image_1_353[47:32]     = Conv_out[462];
    assign  image_1_353[31:16]     = Conv_out[461];
    assign  image_1_353[15:0]      = Conv_out[460];

    assign  image_1_354[143:128]   = Conv_out[521];
    assign  image_1_354[127:112]   = Conv_out[520];
    assign  image_1_354[111:96]    = Conv_out[519];
    assign  image_1_354[95:80]     = Conv_out[491];
    assign  image_1_354[79:64]     = Conv_out[490];
    assign  image_1_354[63:48]     = Conv_out[489];
    assign  image_1_354[47:32]     = Conv_out[461];
    assign  image_1_354[31:16]     = Conv_out[460];
    assign  image_1_354[15:0]      = Conv_out[459];

    assign  image_1_355[143:128]   = Conv_out[520];
    assign  image_1_355[127:112]   = Conv_out[519];
    assign  image_1_355[111:96]    = Conv_out[518];
    assign  image_1_355[95:80]     = Conv_out[490];
    assign  image_1_355[79:64]     = Conv_out[489];
    assign  image_1_355[63:48]     = Conv_out[488];
    assign  image_1_355[47:32]     = Conv_out[460];
    assign  image_1_355[31:16]     = Conv_out[459];
    assign  image_1_355[15:0]      = Conv_out[458];

    assign  image_1_356[143:128]   = Conv_out[519];
    assign  image_1_356[127:112]   = Conv_out[518];
    assign  image_1_356[111:96]    = Conv_out[517];
    assign  image_1_356[95:80]     = Conv_out[489];
    assign  image_1_356[79:64]     = Conv_out[488];
    assign  image_1_356[63:48]     = Conv_out[487];
    assign  image_1_356[47:32]     = Conv_out[459];
    assign  image_1_356[31:16]     = Conv_out[458];
    assign  image_1_356[15:0]      = Conv_out[457];

    assign  image_1_357[143:128]   = Conv_out[518];
    assign  image_1_357[127:112]   = Conv_out[517];
    assign  image_1_357[111:96]    = Conv_out[516];
    assign  image_1_357[95:80]     = Conv_out[488];
    assign  image_1_357[79:64]     = Conv_out[487];
    assign  image_1_357[63:48]     = Conv_out[486];
    assign  image_1_357[47:32]     = Conv_out[458];
    assign  image_1_357[31:16]     = Conv_out[457];
    assign  image_1_357[15:0]      = Conv_out[456];

    assign  image_1_358[143:128]   = Conv_out[517];
    assign  image_1_358[127:112]   = Conv_out[516];
    assign  image_1_358[111:96]    = Conv_out[515];
    assign  image_1_358[95:80]     = Conv_out[487];
    assign  image_1_358[79:64]     = Conv_out[486];
    assign  image_1_358[63:48]     = Conv_out[485];
    assign  image_1_358[47:32]     = Conv_out[457];
    assign  image_1_358[31:16]     = Conv_out[456];
    assign  image_1_358[15:0]      = Conv_out[455];

    assign  image_1_359[143:128]   = Conv_out[516];
    assign  image_1_359[127:112]   = Conv_out[515];
    assign  image_1_359[111:96]    = Conv_out[514];
    assign  image_1_359[95:80]     = Conv_out[486];
    assign  image_1_359[79:64]     = Conv_out[485];
    assign  image_1_359[63:48]     = Conv_out[484];
    assign  image_1_359[47:32]     = Conv_out[456];
    assign  image_1_359[31:16]     = Conv_out[455];
    assign  image_1_359[15:0]      = Conv_out[454];

    assign  image_1_360[143:128]   = Conv_out[515];
    assign  image_1_360[127:112]   = Conv_out[514];
    assign  image_1_360[111:96]    = Conv_out[513];
    assign  image_1_360[95:80]     = Conv_out[485];
    assign  image_1_360[79:64]     = Conv_out[484];
    assign  image_1_360[63:48]     = Conv_out[483];
    assign  image_1_360[47:32]     = Conv_out[455];
    assign  image_1_360[31:16]     = Conv_out[454];
    assign  image_1_360[15:0]      = Conv_out[453];

    assign  image_1_361[143:128]   = Conv_out[514];
    assign  image_1_361[127:112]   = Conv_out[513];
    assign  image_1_361[111:96]    = Conv_out[512];
    assign  image_1_361[95:80]     = Conv_out[484];
    assign  image_1_361[79:64]     = Conv_out[483];
    assign  image_1_361[63:48]     = Conv_out[482];
    assign  image_1_361[47:32]     = Conv_out[454];
    assign  image_1_361[31:16]     = Conv_out[453];
    assign  image_1_361[15:0]      = Conv_out[452];

    assign  image_1_362[143:128]   = Conv_out[513];
    assign  image_1_362[127:112]   = Conv_out[512];
    assign  image_1_362[111:96]    = Conv_out[511];
    assign  image_1_362[95:80]     = Conv_out[483];
    assign  image_1_362[79:64]     = Conv_out[482];
    assign  image_1_362[63:48]     = Conv_out[481];
    assign  image_1_362[47:32]     = Conv_out[453];
    assign  image_1_362[31:16]     = Conv_out[452];
    assign  image_1_362[15:0]      = Conv_out[451];

    assign  image_1_363[143:128]   = Conv_out[512];
    assign  image_1_363[127:112]   = Conv_out[511];
    assign  image_1_363[111:96]    = Conv_out[510];
    assign  image_1_363[95:80]     = Conv_out[482];
    assign  image_1_363[79:64]     = Conv_out[481];
    assign  image_1_363[63:48]     = Conv_out[480];
    assign  image_1_363[47:32]     = Conv_out[452];
    assign  image_1_363[31:16]     = Conv_out[451];
    assign  image_1_363[15:0]      = Conv_out[450];

    assign  image_1_364[143:128]   = Conv_out[509];
    assign  image_1_364[127:112]   = Conv_out[508];
    assign  image_1_364[111:96]    = Conv_out[507];
    assign  image_1_364[95:80]     = Conv_out[479];
    assign  image_1_364[79:64]     = Conv_out[478];
    assign  image_1_364[63:48]     = Conv_out[477];
    assign  image_1_364[47:32]     = Conv_out[449];
    assign  image_1_364[31:16]     = Conv_out[448];
    assign  image_1_364[15:0]      = Conv_out[447];

    assign  image_1_365[143:128]   = Conv_out[508];
    assign  image_1_365[127:112]   = Conv_out[507];
    assign  image_1_365[111:96]    = Conv_out[506];
    assign  image_1_365[95:80]     = Conv_out[478];
    assign  image_1_365[79:64]     = Conv_out[477];
    assign  image_1_365[63:48]     = Conv_out[476];
    assign  image_1_365[47:32]     = Conv_out[448];
    assign  image_1_365[31:16]     = Conv_out[447];
    assign  image_1_365[15:0]      = Conv_out[446];

    assign  image_1_366[143:128]   = Conv_out[507];
    assign  image_1_366[127:112]   = Conv_out[506];
    assign  image_1_366[111:96]    = Conv_out[505];
    assign  image_1_366[95:80]     = Conv_out[477];
    assign  image_1_366[79:64]     = Conv_out[476];
    assign  image_1_366[63:48]     = Conv_out[475];
    assign  image_1_366[47:32]     = Conv_out[447];
    assign  image_1_366[31:16]     = Conv_out[446];
    assign  image_1_366[15:0]      = Conv_out[445];

    assign  image_1_367[143:128]   = Conv_out[506];
    assign  image_1_367[127:112]   = Conv_out[505];
    assign  image_1_367[111:96]    = Conv_out[504];
    assign  image_1_367[95:80]     = Conv_out[476];
    assign  image_1_367[79:64]     = Conv_out[475];
    assign  image_1_367[63:48]     = Conv_out[474];
    assign  image_1_367[47:32]     = Conv_out[446];
    assign  image_1_367[31:16]     = Conv_out[445];
    assign  image_1_367[15:0]      = Conv_out[444];

    assign  image_1_368[143:128]   = Conv_out[505];
    assign  image_1_368[127:112]   = Conv_out[504];
    assign  image_1_368[111:96]    = Conv_out[503];
    assign  image_1_368[95:80]     = Conv_out[475];
    assign  image_1_368[79:64]     = Conv_out[474];
    assign  image_1_368[63:48]     = Conv_out[473];
    assign  image_1_368[47:32]     = Conv_out[445];
    assign  image_1_368[31:16]     = Conv_out[444];
    assign  image_1_368[15:0]      = Conv_out[443];

    assign  image_1_369[143:128]   = Conv_out[504];
    assign  image_1_369[127:112]   = Conv_out[503];
    assign  image_1_369[111:96]    = Conv_out[502];
    assign  image_1_369[95:80]     = Conv_out[474];
    assign  image_1_369[79:64]     = Conv_out[473];
    assign  image_1_369[63:48]     = Conv_out[472];
    assign  image_1_369[47:32]     = Conv_out[444];
    assign  image_1_369[31:16]     = Conv_out[443];
    assign  image_1_369[15:0]      = Conv_out[442];

    assign  image_1_370[143:128]   = Conv_out[503];
    assign  image_1_370[127:112]   = Conv_out[502];
    assign  image_1_370[111:96]    = Conv_out[501];
    assign  image_1_370[95:80]     = Conv_out[473];
    assign  image_1_370[79:64]     = Conv_out[472];
    assign  image_1_370[63:48]     = Conv_out[471];
    assign  image_1_370[47:32]     = Conv_out[443];
    assign  image_1_370[31:16]     = Conv_out[442];
    assign  image_1_370[15:0]      = Conv_out[441];

    assign  image_1_371[143:128]   = Conv_out[502];
    assign  image_1_371[127:112]   = Conv_out[501];
    assign  image_1_371[111:96]    = Conv_out[500];
    assign  image_1_371[95:80]     = Conv_out[472];
    assign  image_1_371[79:64]     = Conv_out[471];
    assign  image_1_371[63:48]     = Conv_out[470];
    assign  image_1_371[47:32]     = Conv_out[442];
    assign  image_1_371[31:16]     = Conv_out[441];
    assign  image_1_371[15:0]      = Conv_out[440];

    assign  image_1_372[143:128]   = Conv_out[501];
    assign  image_1_372[127:112]   = Conv_out[500];
    assign  image_1_372[111:96]    = Conv_out[499];
    assign  image_1_372[95:80]     = Conv_out[471];
    assign  image_1_372[79:64]     = Conv_out[470];
    assign  image_1_372[63:48]     = Conv_out[469];
    assign  image_1_372[47:32]     = Conv_out[441];
    assign  image_1_372[31:16]     = Conv_out[440];
    assign  image_1_372[15:0]      = Conv_out[439];

    assign  image_1_373[143:128]   = Conv_out[500];
    assign  image_1_373[127:112]   = Conv_out[499];
    assign  image_1_373[111:96]    = Conv_out[498];
    assign  image_1_373[95:80]     = Conv_out[470];
    assign  image_1_373[79:64]     = Conv_out[469];
    assign  image_1_373[63:48]     = Conv_out[468];
    assign  image_1_373[47:32]     = Conv_out[440];
    assign  image_1_373[31:16]     = Conv_out[439];
    assign  image_1_373[15:0]      = Conv_out[438];

    assign  image_1_374[143:128]   = Conv_out[499];
    assign  image_1_374[127:112]   = Conv_out[498];
    assign  image_1_374[111:96]    = Conv_out[497];
    assign  image_1_374[95:80]     = Conv_out[469];
    assign  image_1_374[79:64]     = Conv_out[468];
    assign  image_1_374[63:48]     = Conv_out[467];
    assign  image_1_374[47:32]     = Conv_out[439];
    assign  image_1_374[31:16]     = Conv_out[438];
    assign  image_1_374[15:0]      = Conv_out[437];

    assign  image_1_375[143:128]   = Conv_out[498];
    assign  image_1_375[127:112]   = Conv_out[497];
    assign  image_1_375[111:96]    = Conv_out[496];
    assign  image_1_375[95:80]     = Conv_out[468];
    assign  image_1_375[79:64]     = Conv_out[467];
    assign  image_1_375[63:48]     = Conv_out[466];
    assign  image_1_375[47:32]     = Conv_out[438];
    assign  image_1_375[31:16]     = Conv_out[437];
    assign  image_1_375[15:0]      = Conv_out[436];

    assign  image_1_376[143:128]   = Conv_out[497];
    assign  image_1_376[127:112]   = Conv_out[496];
    assign  image_1_376[111:96]    = Conv_out[495];
    assign  image_1_376[95:80]     = Conv_out[467];
    assign  image_1_376[79:64]     = Conv_out[466];
    assign  image_1_376[63:48]     = Conv_out[465];
    assign  image_1_376[47:32]     = Conv_out[437];
    assign  image_1_376[31:16]     = Conv_out[436];
    assign  image_1_376[15:0]      = Conv_out[435];

    assign  image_1_377[143:128]   = Conv_out[496];
    assign  image_1_377[127:112]   = Conv_out[495];
    assign  image_1_377[111:96]    = Conv_out[494];
    assign  image_1_377[95:80]     = Conv_out[466];
    assign  image_1_377[79:64]     = Conv_out[465];
    assign  image_1_377[63:48]     = Conv_out[464];
    assign  image_1_377[47:32]     = Conv_out[436];
    assign  image_1_377[31:16]     = Conv_out[435];
    assign  image_1_377[15:0]      = Conv_out[434];

    assign  image_1_378[143:128]   = Conv_out[495];
    assign  image_1_378[127:112]   = Conv_out[494];
    assign  image_1_378[111:96]    = Conv_out[493];
    assign  image_1_378[95:80]     = Conv_out[465];
    assign  image_1_378[79:64]     = Conv_out[464];
    assign  image_1_378[63:48]     = Conv_out[463];
    assign  image_1_378[47:32]     = Conv_out[435];
    assign  image_1_378[31:16]     = Conv_out[434];
    assign  image_1_378[15:0]      = Conv_out[433];

    assign  image_1_379[143:128]   = Conv_out[494];
    assign  image_1_379[127:112]   = Conv_out[493];
    assign  image_1_379[111:96]    = Conv_out[492];
    assign  image_1_379[95:80]     = Conv_out[464];
    assign  image_1_379[79:64]     = Conv_out[463];
    assign  image_1_379[63:48]     = Conv_out[462];
    assign  image_1_379[47:32]     = Conv_out[434];
    assign  image_1_379[31:16]     = Conv_out[433];
    assign  image_1_379[15:0]      = Conv_out[432];

    assign  image_1_380[143:128]   = Conv_out[493];
    assign  image_1_380[127:112]   = Conv_out[492];
    assign  image_1_380[111:96]    = Conv_out[491];
    assign  image_1_380[95:80]     = Conv_out[463];
    assign  image_1_380[79:64]     = Conv_out[462];
    assign  image_1_380[63:48]     = Conv_out[461];
    assign  image_1_380[47:32]     = Conv_out[433];
    assign  image_1_380[31:16]     = Conv_out[432];
    assign  image_1_380[15:0]      = Conv_out[431];

    assign  image_1_381[143:128]   = Conv_out[492];
    assign  image_1_381[127:112]   = Conv_out[491];
    assign  image_1_381[111:96]    = Conv_out[490];
    assign  image_1_381[95:80]     = Conv_out[462];
    assign  image_1_381[79:64]     = Conv_out[461];
    assign  image_1_381[63:48]     = Conv_out[460];
    assign  image_1_381[47:32]     = Conv_out[432];
    assign  image_1_381[31:16]     = Conv_out[431];
    assign  image_1_381[15:0]      = Conv_out[430];

    assign  image_1_382[143:128]   = Conv_out[491];
    assign  image_1_382[127:112]   = Conv_out[490];
    assign  image_1_382[111:96]    = Conv_out[489];
    assign  image_1_382[95:80]     = Conv_out[461];
    assign  image_1_382[79:64]     = Conv_out[460];
    assign  image_1_382[63:48]     = Conv_out[459];
    assign  image_1_382[47:32]     = Conv_out[431];
    assign  image_1_382[31:16]     = Conv_out[430];
    assign  image_1_382[15:0]      = Conv_out[429];

    assign  image_1_383[143:128]   = Conv_out[490];
    assign  image_1_383[127:112]   = Conv_out[489];
    assign  image_1_383[111:96]    = Conv_out[488];
    assign  image_1_383[95:80]     = Conv_out[460];
    assign  image_1_383[79:64]     = Conv_out[459];
    assign  image_1_383[63:48]     = Conv_out[458];
    assign  image_1_383[47:32]     = Conv_out[430];
    assign  image_1_383[31:16]     = Conv_out[429];
    assign  image_1_383[15:0]      = Conv_out[428];

    assign  image_1_384[143:128]   = Conv_out[489];
    assign  image_1_384[127:112]   = Conv_out[488];
    assign  image_1_384[111:96]    = Conv_out[487];
    assign  image_1_384[95:80]     = Conv_out[459];
    assign  image_1_384[79:64]     = Conv_out[458];
    assign  image_1_384[63:48]     = Conv_out[457];
    assign  image_1_384[47:32]     = Conv_out[429];
    assign  image_1_384[31:16]     = Conv_out[428];
    assign  image_1_384[15:0]      = Conv_out[427];

    assign  image_1_385[143:128]   = Conv_out[488];
    assign  image_1_385[127:112]   = Conv_out[487];
    assign  image_1_385[111:96]    = Conv_out[486];
    assign  image_1_385[95:80]     = Conv_out[458];
    assign  image_1_385[79:64]     = Conv_out[457];
    assign  image_1_385[63:48]     = Conv_out[456];
    assign  image_1_385[47:32]     = Conv_out[428];
    assign  image_1_385[31:16]     = Conv_out[427];
    assign  image_1_385[15:0]      = Conv_out[426];

    assign  image_1_386[143:128]   = Conv_out[487];
    assign  image_1_386[127:112]   = Conv_out[486];
    assign  image_1_386[111:96]    = Conv_out[485];
    assign  image_1_386[95:80]     = Conv_out[457];
    assign  image_1_386[79:64]     = Conv_out[456];
    assign  image_1_386[63:48]     = Conv_out[455];
    assign  image_1_386[47:32]     = Conv_out[427];
    assign  image_1_386[31:16]     = Conv_out[426];
    assign  image_1_386[15:0]      = Conv_out[425];

    assign  image_1_387[143:128]   = Conv_out[486];
    assign  image_1_387[127:112]   = Conv_out[485];
    assign  image_1_387[111:96]    = Conv_out[484];
    assign  image_1_387[95:80]     = Conv_out[456];
    assign  image_1_387[79:64]     = Conv_out[455];
    assign  image_1_387[63:48]     = Conv_out[454];
    assign  image_1_387[47:32]     = Conv_out[426];
    assign  image_1_387[31:16]     = Conv_out[425];
    assign  image_1_387[15:0]      = Conv_out[424];

    assign  image_1_388[143:128]   = Conv_out[485];
    assign  image_1_388[127:112]   = Conv_out[484];
    assign  image_1_388[111:96]    = Conv_out[483];
    assign  image_1_388[95:80]     = Conv_out[455];
    assign  image_1_388[79:64]     = Conv_out[454];
    assign  image_1_388[63:48]     = Conv_out[453];
    assign  image_1_388[47:32]     = Conv_out[425];
    assign  image_1_388[31:16]     = Conv_out[424];
    assign  image_1_388[15:0]      = Conv_out[423];

    assign  image_1_389[143:128]   = Conv_out[484];
    assign  image_1_389[127:112]   = Conv_out[483];
    assign  image_1_389[111:96]    = Conv_out[482];
    assign  image_1_389[95:80]     = Conv_out[454];
    assign  image_1_389[79:64]     = Conv_out[453];
    assign  image_1_389[63:48]     = Conv_out[452];
    assign  image_1_389[47:32]     = Conv_out[424];
    assign  image_1_389[31:16]     = Conv_out[423];
    assign  image_1_389[15:0]      = Conv_out[422];

    assign  image_1_390[143:128]   = Conv_out[483];
    assign  image_1_390[127:112]   = Conv_out[482];
    assign  image_1_390[111:96]    = Conv_out[481];
    assign  image_1_390[95:80]     = Conv_out[453];
    assign  image_1_390[79:64]     = Conv_out[452];
    assign  image_1_390[63:48]     = Conv_out[451];
    assign  image_1_390[47:32]     = Conv_out[423];
    assign  image_1_390[31:16]     = Conv_out[422];
    assign  image_1_390[15:0]      = Conv_out[421];

    assign  image_1_391[143:128]   = Conv_out[482];
    assign  image_1_391[127:112]   = Conv_out[481];
    assign  image_1_391[111:96]    = Conv_out[480];
    assign  image_1_391[95:80]     = Conv_out[452];
    assign  image_1_391[79:64]     = Conv_out[451];
    assign  image_1_391[63:48]     = Conv_out[450];
    assign  image_1_391[47:32]     = Conv_out[422];
    assign  image_1_391[31:16]     = Conv_out[421];
    assign  image_1_391[15:0]      = Conv_out[420];

    assign  image_1_392[143:128]   = Conv_out[479];
    assign  image_1_392[127:112]   = Conv_out[478];
    assign  image_1_392[111:96]    = Conv_out[477];
    assign  image_1_392[95:80]     = Conv_out[449];
    assign  image_1_392[79:64]     = Conv_out[448];
    assign  image_1_392[63:48]     = Conv_out[447];
    assign  image_1_392[47:32]     = Conv_out[419];
    assign  image_1_392[31:16]     = Conv_out[418];
    assign  image_1_392[15:0]      = Conv_out[417];

    assign  image_1_393[143:128]   = Conv_out[478];
    assign  image_1_393[127:112]   = Conv_out[477];
    assign  image_1_393[111:96]    = Conv_out[476];
    assign  image_1_393[95:80]     = Conv_out[448];
    assign  image_1_393[79:64]     = Conv_out[447];
    assign  image_1_393[63:48]     = Conv_out[446];
    assign  image_1_393[47:32]     = Conv_out[418];
    assign  image_1_393[31:16]     = Conv_out[417];
    assign  image_1_393[15:0]      = Conv_out[416];

    assign  image_1_394[143:128]   = Conv_out[477];
    assign  image_1_394[127:112]   = Conv_out[476];
    assign  image_1_394[111:96]    = Conv_out[475];
    assign  image_1_394[95:80]     = Conv_out[447];
    assign  image_1_394[79:64]     = Conv_out[446];
    assign  image_1_394[63:48]     = Conv_out[445];
    assign  image_1_394[47:32]     = Conv_out[417];
    assign  image_1_394[31:16]     = Conv_out[416];
    assign  image_1_394[15:0]      = Conv_out[415];

    assign  image_1_395[143:128]   = Conv_out[476];
    assign  image_1_395[127:112]   = Conv_out[475];
    assign  image_1_395[111:96]    = Conv_out[474];
    assign  image_1_395[95:80]     = Conv_out[446];
    assign  image_1_395[79:64]     = Conv_out[445];
    assign  image_1_395[63:48]     = Conv_out[444];
    assign  image_1_395[47:32]     = Conv_out[416];
    assign  image_1_395[31:16]     = Conv_out[415];
    assign  image_1_395[15:0]      = Conv_out[414];

    assign  image_1_396[143:128]   = Conv_out[475];
    assign  image_1_396[127:112]   = Conv_out[474];
    assign  image_1_396[111:96]    = Conv_out[473];
    assign  image_1_396[95:80]     = Conv_out[445];
    assign  image_1_396[79:64]     = Conv_out[444];
    assign  image_1_396[63:48]     = Conv_out[443];
    assign  image_1_396[47:32]     = Conv_out[415];
    assign  image_1_396[31:16]     = Conv_out[414];
    assign  image_1_396[15:0]      = Conv_out[413];

    assign  image_1_397[143:128]   = Conv_out[474];
    assign  image_1_397[127:112]   = Conv_out[473];
    assign  image_1_397[111:96]    = Conv_out[472];
    assign  image_1_397[95:80]     = Conv_out[444];
    assign  image_1_397[79:64]     = Conv_out[443];
    assign  image_1_397[63:48]     = Conv_out[442];
    assign  image_1_397[47:32]     = Conv_out[414];
    assign  image_1_397[31:16]     = Conv_out[413];
    assign  image_1_397[15:0]      = Conv_out[412];

    assign  image_1_398[143:128]   = Conv_out[473];
    assign  image_1_398[127:112]   = Conv_out[472];
    assign  image_1_398[111:96]    = Conv_out[471];
    assign  image_1_398[95:80]     = Conv_out[443];
    assign  image_1_398[79:64]     = Conv_out[442];
    assign  image_1_398[63:48]     = Conv_out[441];
    assign  image_1_398[47:32]     = Conv_out[413];
    assign  image_1_398[31:16]     = Conv_out[412];
    assign  image_1_398[15:0]      = Conv_out[411];

    assign  image_1_399[143:128]   = Conv_out[472];
    assign  image_1_399[127:112]   = Conv_out[471];
    assign  image_1_399[111:96]    = Conv_out[470];
    assign  image_1_399[95:80]     = Conv_out[442];
    assign  image_1_399[79:64]     = Conv_out[441];
    assign  image_1_399[63:48]     = Conv_out[440];
    assign  image_1_399[47:32]     = Conv_out[412];
    assign  image_1_399[31:16]     = Conv_out[411];
    assign  image_1_399[15:0]      = Conv_out[410];

    assign  image_1_400[143:128]   = Conv_out[471];
    assign  image_1_400[127:112]   = Conv_out[470];
    assign  image_1_400[111:96]    = Conv_out[469];
    assign  image_1_400[95:80]     = Conv_out[441];
    assign  image_1_400[79:64]     = Conv_out[440];
    assign  image_1_400[63:48]     = Conv_out[439];
    assign  image_1_400[47:32]     = Conv_out[411];
    assign  image_1_400[31:16]     = Conv_out[410];
    assign  image_1_400[15:0]      = Conv_out[409];

    assign  image_1_401[143:128]   = Conv_out[470];
    assign  image_1_401[127:112]   = Conv_out[469];
    assign  image_1_401[111:96]    = Conv_out[468];
    assign  image_1_401[95:80]     = Conv_out[440];
    assign  image_1_401[79:64]     = Conv_out[439];
    assign  image_1_401[63:48]     = Conv_out[438];
    assign  image_1_401[47:32]     = Conv_out[410];
    assign  image_1_401[31:16]     = Conv_out[409];
    assign  image_1_401[15:0]      = Conv_out[408];

    assign  image_1_402[143:128]   = Conv_out[469];
    assign  image_1_402[127:112]   = Conv_out[468];
    assign  image_1_402[111:96]    = Conv_out[467];
    assign  image_1_402[95:80]     = Conv_out[439];
    assign  image_1_402[79:64]     = Conv_out[438];
    assign  image_1_402[63:48]     = Conv_out[437];
    assign  image_1_402[47:32]     = Conv_out[409];
    assign  image_1_402[31:16]     = Conv_out[408];
    assign  image_1_402[15:0]      = Conv_out[407];

    assign  image_1_403[143:128]   = Conv_out[468];
    assign  image_1_403[127:112]   = Conv_out[467];
    assign  image_1_403[111:96]    = Conv_out[466];
    assign  image_1_403[95:80]     = Conv_out[438];
    assign  image_1_403[79:64]     = Conv_out[437];
    assign  image_1_403[63:48]     = Conv_out[436];
    assign  image_1_403[47:32]     = Conv_out[408];
    assign  image_1_403[31:16]     = Conv_out[407];
    assign  image_1_403[15:0]      = Conv_out[406];

    assign  image_1_404[143:128]   = Conv_out[467];
    assign  image_1_404[127:112]   = Conv_out[466];
    assign  image_1_404[111:96]    = Conv_out[465];
    assign  image_1_404[95:80]     = Conv_out[437];
    assign  image_1_404[79:64]     = Conv_out[436];
    assign  image_1_404[63:48]     = Conv_out[435];
    assign  image_1_404[47:32]     = Conv_out[407];
    assign  image_1_404[31:16]     = Conv_out[406];
    assign  image_1_404[15:0]      = Conv_out[405];

    assign  image_1_405[143:128]   = Conv_out[466];
    assign  image_1_405[127:112]   = Conv_out[465];
    assign  image_1_405[111:96]    = Conv_out[464];
    assign  image_1_405[95:80]     = Conv_out[436];
    assign  image_1_405[79:64]     = Conv_out[435];
    assign  image_1_405[63:48]     = Conv_out[434];
    assign  image_1_405[47:32]     = Conv_out[406];
    assign  image_1_405[31:16]     = Conv_out[405];
    assign  image_1_405[15:0]      = Conv_out[404];

    assign  image_1_406[143:128]   = Conv_out[465];
    assign  image_1_406[127:112]   = Conv_out[464];
    assign  image_1_406[111:96]    = Conv_out[463];
    assign  image_1_406[95:80]     = Conv_out[435];
    assign  image_1_406[79:64]     = Conv_out[434];
    assign  image_1_406[63:48]     = Conv_out[433];
    assign  image_1_406[47:32]     = Conv_out[405];
    assign  image_1_406[31:16]     = Conv_out[404];
    assign  image_1_406[15:0]      = Conv_out[403];

    assign  image_1_407[143:128]   = Conv_out[464];
    assign  image_1_407[127:112]   = Conv_out[463];
    assign  image_1_407[111:96]    = Conv_out[462];
    assign  image_1_407[95:80]     = Conv_out[434];
    assign  image_1_407[79:64]     = Conv_out[433];
    assign  image_1_407[63:48]     = Conv_out[432];
    assign  image_1_407[47:32]     = Conv_out[404];
    assign  image_1_407[31:16]     = Conv_out[403];
    assign  image_1_407[15:0]      = Conv_out[402];

    assign  image_1_408[143:128]   = Conv_out[463];
    assign  image_1_408[127:112]   = Conv_out[462];
    assign  image_1_408[111:96]    = Conv_out[461];
    assign  image_1_408[95:80]     = Conv_out[433];
    assign  image_1_408[79:64]     = Conv_out[432];
    assign  image_1_408[63:48]     = Conv_out[431];
    assign  image_1_408[47:32]     = Conv_out[403];
    assign  image_1_408[31:16]     = Conv_out[402];
    assign  image_1_408[15:0]      = Conv_out[401];

    assign  image_1_409[143:128]   = Conv_out[462];
    assign  image_1_409[127:112]   = Conv_out[461];
    assign  image_1_409[111:96]    = Conv_out[460];
    assign  image_1_409[95:80]     = Conv_out[432];
    assign  image_1_409[79:64]     = Conv_out[431];
    assign  image_1_409[63:48]     = Conv_out[430];
    assign  image_1_409[47:32]     = Conv_out[402];
    assign  image_1_409[31:16]     = Conv_out[401];
    assign  image_1_409[15:0]      = Conv_out[400];

    assign  image_1_410[143:128]   = Conv_out[461];
    assign  image_1_410[127:112]   = Conv_out[460];
    assign  image_1_410[111:96]    = Conv_out[459];
    assign  image_1_410[95:80]     = Conv_out[431];
    assign  image_1_410[79:64]     = Conv_out[430];
    assign  image_1_410[63:48]     = Conv_out[429];
    assign  image_1_410[47:32]     = Conv_out[401];
    assign  image_1_410[31:16]     = Conv_out[400];
    assign  image_1_410[15:0]      = Conv_out[399];

    assign  image_1_411[143:128]   = Conv_out[460];
    assign  image_1_411[127:112]   = Conv_out[459];
    assign  image_1_411[111:96]    = Conv_out[458];
    assign  image_1_411[95:80]     = Conv_out[430];
    assign  image_1_411[79:64]     = Conv_out[429];
    assign  image_1_411[63:48]     = Conv_out[428];
    assign  image_1_411[47:32]     = Conv_out[400];
    assign  image_1_411[31:16]     = Conv_out[399];
    assign  image_1_411[15:0]      = Conv_out[398];

    assign  image_1_412[143:128]   = Conv_out[459];
    assign  image_1_412[127:112]   = Conv_out[458];
    assign  image_1_412[111:96]    = Conv_out[457];
    assign  image_1_412[95:80]     = Conv_out[429];
    assign  image_1_412[79:64]     = Conv_out[428];
    assign  image_1_412[63:48]     = Conv_out[427];
    assign  image_1_412[47:32]     = Conv_out[399];
    assign  image_1_412[31:16]     = Conv_out[398];
    assign  image_1_412[15:0]      = Conv_out[397];

    assign  image_1_413[143:128]   = Conv_out[458];
    assign  image_1_413[127:112]   = Conv_out[457];
    assign  image_1_413[111:96]    = Conv_out[456];
    assign  image_1_413[95:80]     = Conv_out[428];
    assign  image_1_413[79:64]     = Conv_out[427];
    assign  image_1_413[63:48]     = Conv_out[426];
    assign  image_1_413[47:32]     = Conv_out[398];
    assign  image_1_413[31:16]     = Conv_out[397];
    assign  image_1_413[15:0]      = Conv_out[396];

    assign  image_1_414[143:128]   = Conv_out[457];
    assign  image_1_414[127:112]   = Conv_out[456];
    assign  image_1_414[111:96]    = Conv_out[455];
    assign  image_1_414[95:80]     = Conv_out[427];
    assign  image_1_414[79:64]     = Conv_out[426];
    assign  image_1_414[63:48]     = Conv_out[425];
    assign  image_1_414[47:32]     = Conv_out[397];
    assign  image_1_414[31:16]     = Conv_out[396];
    assign  image_1_414[15:0]      = Conv_out[395];

    assign  image_1_415[143:128]   = Conv_out[456];
    assign  image_1_415[127:112]   = Conv_out[455];
    assign  image_1_415[111:96]    = Conv_out[454];
    assign  image_1_415[95:80]     = Conv_out[426];
    assign  image_1_415[79:64]     = Conv_out[425];
    assign  image_1_415[63:48]     = Conv_out[424];
    assign  image_1_415[47:32]     = Conv_out[396];
    assign  image_1_415[31:16]     = Conv_out[395];
    assign  image_1_415[15:0]      = Conv_out[394];

    assign  image_1_416[143:128]   = Conv_out[455];
    assign  image_1_416[127:112]   = Conv_out[454];
    assign  image_1_416[111:96]    = Conv_out[453];
    assign  image_1_416[95:80]     = Conv_out[425];
    assign  image_1_416[79:64]     = Conv_out[424];
    assign  image_1_416[63:48]     = Conv_out[423];
    assign  image_1_416[47:32]     = Conv_out[395];
    assign  image_1_416[31:16]     = Conv_out[394];
    assign  image_1_416[15:0]      = Conv_out[393];

    assign  image_1_417[143:128]   = Conv_out[454];
    assign  image_1_417[127:112]   = Conv_out[453];
    assign  image_1_417[111:96]    = Conv_out[452];
    assign  image_1_417[95:80]     = Conv_out[424];
    assign  image_1_417[79:64]     = Conv_out[423];
    assign  image_1_417[63:48]     = Conv_out[422];
    assign  image_1_417[47:32]     = Conv_out[394];
    assign  image_1_417[31:16]     = Conv_out[393];
    assign  image_1_417[15:0]      = Conv_out[392];

    assign  image_1_418[143:128]   = Conv_out[453];
    assign  image_1_418[127:112]   = Conv_out[452];
    assign  image_1_418[111:96]    = Conv_out[451];
    assign  image_1_418[95:80]     = Conv_out[423];
    assign  image_1_418[79:64]     = Conv_out[422];
    assign  image_1_418[63:48]     = Conv_out[421];
    assign  image_1_418[47:32]     = Conv_out[393];
    assign  image_1_418[31:16]     = Conv_out[392];
    assign  image_1_418[15:0]      = Conv_out[391];

    assign  image_1_419[143:128]   = Conv_out[452];
    assign  image_1_419[127:112]   = Conv_out[451];
    assign  image_1_419[111:96]    = Conv_out[450];
    assign  image_1_419[95:80]     = Conv_out[422];
    assign  image_1_419[79:64]     = Conv_out[421];
    assign  image_1_419[63:48]     = Conv_out[420];
    assign  image_1_419[47:32]     = Conv_out[392];
    assign  image_1_419[31:16]     = Conv_out[391];
    assign  image_1_419[15:0]      = Conv_out[390];

    assign  image_1_420[143:128]   = Conv_out[449];
    assign  image_1_420[127:112]   = Conv_out[448];
    assign  image_1_420[111:96]    = Conv_out[447];
    assign  image_1_420[95:80]     = Conv_out[419];
    assign  image_1_420[79:64]     = Conv_out[418];
    assign  image_1_420[63:48]     = Conv_out[417];
    assign  image_1_420[47:32]     = Conv_out[389];
    assign  image_1_420[31:16]     = Conv_out[388];
    assign  image_1_420[15:0]      = Conv_out[387];

    assign  image_1_421[143:128]   = Conv_out[448];
    assign  image_1_421[127:112]   = Conv_out[447];
    assign  image_1_421[111:96]    = Conv_out[446];
    assign  image_1_421[95:80]     = Conv_out[418];
    assign  image_1_421[79:64]     = Conv_out[417];
    assign  image_1_421[63:48]     = Conv_out[416];
    assign  image_1_421[47:32]     = Conv_out[388];
    assign  image_1_421[31:16]     = Conv_out[387];
    assign  image_1_421[15:0]      = Conv_out[386];

    assign  image_1_422[143:128]   = Conv_out[447];
    assign  image_1_422[127:112]   = Conv_out[446];
    assign  image_1_422[111:96]    = Conv_out[445];
    assign  image_1_422[95:80]     = Conv_out[417];
    assign  image_1_422[79:64]     = Conv_out[416];
    assign  image_1_422[63:48]     = Conv_out[415];
    assign  image_1_422[47:32]     = Conv_out[387];
    assign  image_1_422[31:16]     = Conv_out[386];
    assign  image_1_422[15:0]      = Conv_out[385];

    assign  image_1_423[143:128]   = Conv_out[446];
    assign  image_1_423[127:112]   = Conv_out[445];
    assign  image_1_423[111:96]    = Conv_out[444];
    assign  image_1_423[95:80]     = Conv_out[416];
    assign  image_1_423[79:64]     = Conv_out[415];
    assign  image_1_423[63:48]     = Conv_out[414];
    assign  image_1_423[47:32]     = Conv_out[386];
    assign  image_1_423[31:16]     = Conv_out[385];
    assign  image_1_423[15:0]      = Conv_out[384];

    assign  image_1_424[143:128]   = Conv_out[445];
    assign  image_1_424[127:112]   = Conv_out[444];
    assign  image_1_424[111:96]    = Conv_out[443];
    assign  image_1_424[95:80]     = Conv_out[415];
    assign  image_1_424[79:64]     = Conv_out[414];
    assign  image_1_424[63:48]     = Conv_out[413];
    assign  image_1_424[47:32]     = Conv_out[385];
    assign  image_1_424[31:16]     = Conv_out[384];
    assign  image_1_424[15:0]      = Conv_out[383];

    assign  image_1_425[143:128]   = Conv_out[444];
    assign  image_1_425[127:112]   = Conv_out[443];
    assign  image_1_425[111:96]    = Conv_out[442];
    assign  image_1_425[95:80]     = Conv_out[414];
    assign  image_1_425[79:64]     = Conv_out[413];
    assign  image_1_425[63:48]     = Conv_out[412];
    assign  image_1_425[47:32]     = Conv_out[384];
    assign  image_1_425[31:16]     = Conv_out[383];
    assign  image_1_425[15:0]      = Conv_out[382];

    assign  image_1_426[143:128]   = Conv_out[443];
    assign  image_1_426[127:112]   = Conv_out[442];
    assign  image_1_426[111:96]    = Conv_out[441];
    assign  image_1_426[95:80]     = Conv_out[413];
    assign  image_1_426[79:64]     = Conv_out[412];
    assign  image_1_426[63:48]     = Conv_out[411];
    assign  image_1_426[47:32]     = Conv_out[383];
    assign  image_1_426[31:16]     = Conv_out[382];
    assign  image_1_426[15:0]      = Conv_out[381];

    assign  image_1_427[143:128]   = Conv_out[442];
    assign  image_1_427[127:112]   = Conv_out[441];
    assign  image_1_427[111:96]    = Conv_out[440];
    assign  image_1_427[95:80]     = Conv_out[412];
    assign  image_1_427[79:64]     = Conv_out[411];
    assign  image_1_427[63:48]     = Conv_out[410];
    assign  image_1_427[47:32]     = Conv_out[382];
    assign  image_1_427[31:16]     = Conv_out[381];
    assign  image_1_427[15:0]      = Conv_out[380];

    assign  image_1_428[143:128]   = Conv_out[441];
    assign  image_1_428[127:112]   = Conv_out[440];
    assign  image_1_428[111:96]    = Conv_out[439];
    assign  image_1_428[95:80]     = Conv_out[411];
    assign  image_1_428[79:64]     = Conv_out[410];
    assign  image_1_428[63:48]     = Conv_out[409];
    assign  image_1_428[47:32]     = Conv_out[381];
    assign  image_1_428[31:16]     = Conv_out[380];
    assign  image_1_428[15:0]      = Conv_out[379];

    assign  image_1_429[143:128]   = Conv_out[440];
    assign  image_1_429[127:112]   = Conv_out[439];
    assign  image_1_429[111:96]    = Conv_out[438];
    assign  image_1_429[95:80]     = Conv_out[410];
    assign  image_1_429[79:64]     = Conv_out[409];
    assign  image_1_429[63:48]     = Conv_out[408];
    assign  image_1_429[47:32]     = Conv_out[380];
    assign  image_1_429[31:16]     = Conv_out[379];
    assign  image_1_429[15:0]      = Conv_out[378];

    assign  image_1_430[143:128]   = Conv_out[439];
    assign  image_1_430[127:112]   = Conv_out[438];
    assign  image_1_430[111:96]    = Conv_out[437];
    assign  image_1_430[95:80]     = Conv_out[409];
    assign  image_1_430[79:64]     = Conv_out[408];
    assign  image_1_430[63:48]     = Conv_out[407];
    assign  image_1_430[47:32]     = Conv_out[379];
    assign  image_1_430[31:16]     = Conv_out[378];
    assign  image_1_430[15:0]      = Conv_out[377];

    assign  image_1_431[143:128]   = Conv_out[438];
    assign  image_1_431[127:112]   = Conv_out[437];
    assign  image_1_431[111:96]    = Conv_out[436];
    assign  image_1_431[95:80]     = Conv_out[408];
    assign  image_1_431[79:64]     = Conv_out[407];
    assign  image_1_431[63:48]     = Conv_out[406];
    assign  image_1_431[47:32]     = Conv_out[378];
    assign  image_1_431[31:16]     = Conv_out[377];
    assign  image_1_431[15:0]      = Conv_out[376];

    assign  image_1_432[143:128]   = Conv_out[437];
    assign  image_1_432[127:112]   = Conv_out[436];
    assign  image_1_432[111:96]    = Conv_out[435];
    assign  image_1_432[95:80]     = Conv_out[407];
    assign  image_1_432[79:64]     = Conv_out[406];
    assign  image_1_432[63:48]     = Conv_out[405];
    assign  image_1_432[47:32]     = Conv_out[377];
    assign  image_1_432[31:16]     = Conv_out[376];
    assign  image_1_432[15:0]      = Conv_out[375];

    assign  image_1_433[143:128]   = Conv_out[436];
    assign  image_1_433[127:112]   = Conv_out[435];
    assign  image_1_433[111:96]    = Conv_out[434];
    assign  image_1_433[95:80]     = Conv_out[406];
    assign  image_1_433[79:64]     = Conv_out[405];
    assign  image_1_433[63:48]     = Conv_out[404];
    assign  image_1_433[47:32]     = Conv_out[376];
    assign  image_1_433[31:16]     = Conv_out[375];
    assign  image_1_433[15:0]      = Conv_out[374];

    assign  image_1_434[143:128]   = Conv_out[435];
    assign  image_1_434[127:112]   = Conv_out[434];
    assign  image_1_434[111:96]    = Conv_out[433];
    assign  image_1_434[95:80]     = Conv_out[405];
    assign  image_1_434[79:64]     = Conv_out[404];
    assign  image_1_434[63:48]     = Conv_out[403];
    assign  image_1_434[47:32]     = Conv_out[375];
    assign  image_1_434[31:16]     = Conv_out[374];
    assign  image_1_434[15:0]      = Conv_out[373];

    assign  image_1_435[143:128]   = Conv_out[434];
    assign  image_1_435[127:112]   = Conv_out[433];
    assign  image_1_435[111:96]    = Conv_out[432];
    assign  image_1_435[95:80]     = Conv_out[404];
    assign  image_1_435[79:64]     = Conv_out[403];
    assign  image_1_435[63:48]     = Conv_out[402];
    assign  image_1_435[47:32]     = Conv_out[374];
    assign  image_1_435[31:16]     = Conv_out[373];
    assign  image_1_435[15:0]      = Conv_out[372];

    assign  image_1_436[143:128]   = Conv_out[433];
    assign  image_1_436[127:112]   = Conv_out[432];
    assign  image_1_436[111:96]    = Conv_out[431];
    assign  image_1_436[95:80]     = Conv_out[403];
    assign  image_1_436[79:64]     = Conv_out[402];
    assign  image_1_436[63:48]     = Conv_out[401];
    assign  image_1_436[47:32]     = Conv_out[373];
    assign  image_1_436[31:16]     = Conv_out[372];
    assign  image_1_436[15:0]      = Conv_out[371];

    assign  image_1_437[143:128]   = Conv_out[432];
    assign  image_1_437[127:112]   = Conv_out[431];
    assign  image_1_437[111:96]    = Conv_out[430];
    assign  image_1_437[95:80]     = Conv_out[402];
    assign  image_1_437[79:64]     = Conv_out[401];
    assign  image_1_437[63:48]     = Conv_out[400];
    assign  image_1_437[47:32]     = Conv_out[372];
    assign  image_1_437[31:16]     = Conv_out[371];
    assign  image_1_437[15:0]      = Conv_out[370];

    assign  image_1_438[143:128]   = Conv_out[431];
    assign  image_1_438[127:112]   = Conv_out[430];
    assign  image_1_438[111:96]    = Conv_out[429];
    assign  image_1_438[95:80]     = Conv_out[401];
    assign  image_1_438[79:64]     = Conv_out[400];
    assign  image_1_438[63:48]     = Conv_out[399];
    assign  image_1_438[47:32]     = Conv_out[371];
    assign  image_1_438[31:16]     = Conv_out[370];
    assign  image_1_438[15:0]      = Conv_out[369];

    assign  image_1_439[143:128]   = Conv_out[430];
    assign  image_1_439[127:112]   = Conv_out[429];
    assign  image_1_439[111:96]    = Conv_out[428];
    assign  image_1_439[95:80]     = Conv_out[400];
    assign  image_1_439[79:64]     = Conv_out[399];
    assign  image_1_439[63:48]     = Conv_out[398];
    assign  image_1_439[47:32]     = Conv_out[370];
    assign  image_1_439[31:16]     = Conv_out[369];
    assign  image_1_439[15:0]      = Conv_out[368];

    assign  image_1_440[143:128]   = Conv_out[429];
    assign  image_1_440[127:112]   = Conv_out[428];
    assign  image_1_440[111:96]    = Conv_out[427];
    assign  image_1_440[95:80]     = Conv_out[399];
    assign  image_1_440[79:64]     = Conv_out[398];
    assign  image_1_440[63:48]     = Conv_out[397];
    assign  image_1_440[47:32]     = Conv_out[369];
    assign  image_1_440[31:16]     = Conv_out[368];
    assign  image_1_440[15:0]      = Conv_out[367];

    assign  image_1_441[143:128]   = Conv_out[428];
    assign  image_1_441[127:112]   = Conv_out[427];
    assign  image_1_441[111:96]    = Conv_out[426];
    assign  image_1_441[95:80]     = Conv_out[398];
    assign  image_1_441[79:64]     = Conv_out[397];
    assign  image_1_441[63:48]     = Conv_out[396];
    assign  image_1_441[47:32]     = Conv_out[368];
    assign  image_1_441[31:16]     = Conv_out[367];
    assign  image_1_441[15:0]      = Conv_out[366];

    assign  image_1_442[143:128]   = Conv_out[427];
    assign  image_1_442[127:112]   = Conv_out[426];
    assign  image_1_442[111:96]    = Conv_out[425];
    assign  image_1_442[95:80]     = Conv_out[397];
    assign  image_1_442[79:64]     = Conv_out[396];
    assign  image_1_442[63:48]     = Conv_out[395];
    assign  image_1_442[47:32]     = Conv_out[367];
    assign  image_1_442[31:16]     = Conv_out[366];
    assign  image_1_442[15:0]      = Conv_out[365];

    assign  image_1_443[143:128]   = Conv_out[426];
    assign  image_1_443[127:112]   = Conv_out[425];
    assign  image_1_443[111:96]    = Conv_out[424];
    assign  image_1_443[95:80]     = Conv_out[396];
    assign  image_1_443[79:64]     = Conv_out[395];
    assign  image_1_443[63:48]     = Conv_out[394];
    assign  image_1_443[47:32]     = Conv_out[366];
    assign  image_1_443[31:16]     = Conv_out[365];
    assign  image_1_443[15:0]      = Conv_out[364];

    assign  image_1_444[143:128]   = Conv_out[425];
    assign  image_1_444[127:112]   = Conv_out[424];
    assign  image_1_444[111:96]    = Conv_out[423];
    assign  image_1_444[95:80]     = Conv_out[395];
    assign  image_1_444[79:64]     = Conv_out[394];
    assign  image_1_444[63:48]     = Conv_out[393];
    assign  image_1_444[47:32]     = Conv_out[365];
    assign  image_1_444[31:16]     = Conv_out[364];
    assign  image_1_444[15:0]      = Conv_out[363];

    assign  image_1_445[143:128]   = Conv_out[424];
    assign  image_1_445[127:112]   = Conv_out[423];
    assign  image_1_445[111:96]    = Conv_out[422];
    assign  image_1_445[95:80]     = Conv_out[394];
    assign  image_1_445[79:64]     = Conv_out[393];
    assign  image_1_445[63:48]     = Conv_out[392];
    assign  image_1_445[47:32]     = Conv_out[364];
    assign  image_1_445[31:16]     = Conv_out[363];
    assign  image_1_445[15:0]      = Conv_out[362];

    assign  image_1_446[143:128]   = Conv_out[423];
    assign  image_1_446[127:112]   = Conv_out[422];
    assign  image_1_446[111:96]    = Conv_out[421];
    assign  image_1_446[95:80]     = Conv_out[393];
    assign  image_1_446[79:64]     = Conv_out[392];
    assign  image_1_446[63:48]     = Conv_out[391];
    assign  image_1_446[47:32]     = Conv_out[363];
    assign  image_1_446[31:16]     = Conv_out[362];
    assign  image_1_446[15:0]      = Conv_out[361];

    assign  image_1_447[143:128]   = Conv_out[422];
    assign  image_1_447[127:112]   = Conv_out[421];
    assign  image_1_447[111:96]    = Conv_out[420];
    assign  image_1_447[95:80]     = Conv_out[392];
    assign  image_1_447[79:64]     = Conv_out[391];
    assign  image_1_447[63:48]     = Conv_out[390];
    assign  image_1_447[47:32]     = Conv_out[362];
    assign  image_1_447[31:16]     = Conv_out[361];
    assign  image_1_447[15:0]      = Conv_out[360];

    assign  image_1_448[143:128]   = Conv_out[419];
    assign  image_1_448[127:112]   = Conv_out[418];
    assign  image_1_448[111:96]    = Conv_out[417];
    assign  image_1_448[95:80]     = Conv_out[389];
    assign  image_1_448[79:64]     = Conv_out[388];
    assign  image_1_448[63:48]     = Conv_out[387];
    assign  image_1_448[47:32]     = Conv_out[359];
    assign  image_1_448[31:16]     = Conv_out[358];
    assign  image_1_448[15:0]      = Conv_out[357];

    assign  image_1_449[143:128]   = Conv_out[418];
    assign  image_1_449[127:112]   = Conv_out[417];
    assign  image_1_449[111:96]    = Conv_out[416];
    assign  image_1_449[95:80]     = Conv_out[388];
    assign  image_1_449[79:64]     = Conv_out[387];
    assign  image_1_449[63:48]     = Conv_out[386];
    assign  image_1_449[47:32]     = Conv_out[358];
    assign  image_1_449[31:16]     = Conv_out[357];
    assign  image_1_449[15:0]      = Conv_out[356];

    assign  image_1_450[143:128]   = Conv_out[417];
    assign  image_1_450[127:112]   = Conv_out[416];
    assign  image_1_450[111:96]    = Conv_out[415];
    assign  image_1_450[95:80]     = Conv_out[387];
    assign  image_1_450[79:64]     = Conv_out[386];
    assign  image_1_450[63:48]     = Conv_out[385];
    assign  image_1_450[47:32]     = Conv_out[357];
    assign  image_1_450[31:16]     = Conv_out[356];
    assign  image_1_450[15:0]      = Conv_out[355];

    assign  image_1_451[143:128]   = Conv_out[416];
    assign  image_1_451[127:112]   = Conv_out[415];
    assign  image_1_451[111:96]    = Conv_out[414];
    assign  image_1_451[95:80]     = Conv_out[386];
    assign  image_1_451[79:64]     = Conv_out[385];
    assign  image_1_451[63:48]     = Conv_out[384];
    assign  image_1_451[47:32]     = Conv_out[356];
    assign  image_1_451[31:16]     = Conv_out[355];
    assign  image_1_451[15:0]      = Conv_out[354];

    assign  image_1_452[143:128]   = Conv_out[415];
    assign  image_1_452[127:112]   = Conv_out[414];
    assign  image_1_452[111:96]    = Conv_out[413];
    assign  image_1_452[95:80]     = Conv_out[385];
    assign  image_1_452[79:64]     = Conv_out[384];
    assign  image_1_452[63:48]     = Conv_out[383];
    assign  image_1_452[47:32]     = Conv_out[355];
    assign  image_1_452[31:16]     = Conv_out[354];
    assign  image_1_452[15:0]      = Conv_out[353];

    assign  image_1_453[143:128]   = Conv_out[414];
    assign  image_1_453[127:112]   = Conv_out[413];
    assign  image_1_453[111:96]    = Conv_out[412];
    assign  image_1_453[95:80]     = Conv_out[384];
    assign  image_1_453[79:64]     = Conv_out[383];
    assign  image_1_453[63:48]     = Conv_out[382];
    assign  image_1_453[47:32]     = Conv_out[354];
    assign  image_1_453[31:16]     = Conv_out[353];
    assign  image_1_453[15:0]      = Conv_out[352];

    assign  image_1_454[143:128]   = Conv_out[413];
    assign  image_1_454[127:112]   = Conv_out[412];
    assign  image_1_454[111:96]    = Conv_out[411];
    assign  image_1_454[95:80]     = Conv_out[383];
    assign  image_1_454[79:64]     = Conv_out[382];
    assign  image_1_454[63:48]     = Conv_out[381];
    assign  image_1_454[47:32]     = Conv_out[353];
    assign  image_1_454[31:16]     = Conv_out[352];
    assign  image_1_454[15:0]      = Conv_out[351];

    assign  image_1_455[143:128]   = Conv_out[412];
    assign  image_1_455[127:112]   = Conv_out[411];
    assign  image_1_455[111:96]    = Conv_out[410];
    assign  image_1_455[95:80]     = Conv_out[382];
    assign  image_1_455[79:64]     = Conv_out[381];
    assign  image_1_455[63:48]     = Conv_out[380];
    assign  image_1_455[47:32]     = Conv_out[352];
    assign  image_1_455[31:16]     = Conv_out[351];
    assign  image_1_455[15:0]      = Conv_out[350];

    assign  image_1_456[143:128]   = Conv_out[411];
    assign  image_1_456[127:112]   = Conv_out[410];
    assign  image_1_456[111:96]    = Conv_out[409];
    assign  image_1_456[95:80]     = Conv_out[381];
    assign  image_1_456[79:64]     = Conv_out[380];
    assign  image_1_456[63:48]     = Conv_out[379];
    assign  image_1_456[47:32]     = Conv_out[351];
    assign  image_1_456[31:16]     = Conv_out[350];
    assign  image_1_456[15:0]      = Conv_out[349];

    assign  image_1_457[143:128]   = Conv_out[410];
    assign  image_1_457[127:112]   = Conv_out[409];
    assign  image_1_457[111:96]    = Conv_out[408];
    assign  image_1_457[95:80]     = Conv_out[380];
    assign  image_1_457[79:64]     = Conv_out[379];
    assign  image_1_457[63:48]     = Conv_out[378];
    assign  image_1_457[47:32]     = Conv_out[350];
    assign  image_1_457[31:16]     = Conv_out[349];
    assign  image_1_457[15:0]      = Conv_out[348];

    assign  image_1_458[143:128]   = Conv_out[409];
    assign  image_1_458[127:112]   = Conv_out[408];
    assign  image_1_458[111:96]    = Conv_out[407];
    assign  image_1_458[95:80]     = Conv_out[379];
    assign  image_1_458[79:64]     = Conv_out[378];
    assign  image_1_458[63:48]     = Conv_out[377];
    assign  image_1_458[47:32]     = Conv_out[349];
    assign  image_1_458[31:16]     = Conv_out[348];
    assign  image_1_458[15:0]      = Conv_out[347];

    assign  image_1_459[143:128]   = Conv_out[408];
    assign  image_1_459[127:112]   = Conv_out[407];
    assign  image_1_459[111:96]    = Conv_out[406];
    assign  image_1_459[95:80]     = Conv_out[378];
    assign  image_1_459[79:64]     = Conv_out[377];
    assign  image_1_459[63:48]     = Conv_out[376];
    assign  image_1_459[47:32]     = Conv_out[348];
    assign  image_1_459[31:16]     = Conv_out[347];
    assign  image_1_459[15:0]      = Conv_out[346];

    assign  image_1_460[143:128]   = Conv_out[407];
    assign  image_1_460[127:112]   = Conv_out[406];
    assign  image_1_460[111:96]    = Conv_out[405];
    assign  image_1_460[95:80]     = Conv_out[377];
    assign  image_1_460[79:64]     = Conv_out[376];
    assign  image_1_460[63:48]     = Conv_out[375];
    assign  image_1_460[47:32]     = Conv_out[347];
    assign  image_1_460[31:16]     = Conv_out[346];
    assign  image_1_460[15:0]      = Conv_out[345];

    assign  image_1_461[143:128]   = Conv_out[406];
    assign  image_1_461[127:112]   = Conv_out[405];
    assign  image_1_461[111:96]    = Conv_out[404];
    assign  image_1_461[95:80]     = Conv_out[376];
    assign  image_1_461[79:64]     = Conv_out[375];
    assign  image_1_461[63:48]     = Conv_out[374];
    assign  image_1_461[47:32]     = Conv_out[346];
    assign  image_1_461[31:16]     = Conv_out[345];
    assign  image_1_461[15:0]      = Conv_out[344];

    assign  image_1_462[143:128]   = Conv_out[405];
    assign  image_1_462[127:112]   = Conv_out[404];
    assign  image_1_462[111:96]    = Conv_out[403];
    assign  image_1_462[95:80]     = Conv_out[375];
    assign  image_1_462[79:64]     = Conv_out[374];
    assign  image_1_462[63:48]     = Conv_out[373];
    assign  image_1_462[47:32]     = Conv_out[345];
    assign  image_1_462[31:16]     = Conv_out[344];
    assign  image_1_462[15:0]      = Conv_out[343];

    assign  image_1_463[143:128]   = Conv_out[404];
    assign  image_1_463[127:112]   = Conv_out[403];
    assign  image_1_463[111:96]    = Conv_out[402];
    assign  image_1_463[95:80]     = Conv_out[374];
    assign  image_1_463[79:64]     = Conv_out[373];
    assign  image_1_463[63:48]     = Conv_out[372];
    assign  image_1_463[47:32]     = Conv_out[344];
    assign  image_1_463[31:16]     = Conv_out[343];
    assign  image_1_463[15:0]      = Conv_out[342];

    assign  image_1_464[143:128]   = Conv_out[403];
    assign  image_1_464[127:112]   = Conv_out[402];
    assign  image_1_464[111:96]    = Conv_out[401];
    assign  image_1_464[95:80]     = Conv_out[373];
    assign  image_1_464[79:64]     = Conv_out[372];
    assign  image_1_464[63:48]     = Conv_out[371];
    assign  image_1_464[47:32]     = Conv_out[343];
    assign  image_1_464[31:16]     = Conv_out[342];
    assign  image_1_464[15:0]      = Conv_out[341];

    assign  image_1_465[143:128]   = Conv_out[402];
    assign  image_1_465[127:112]   = Conv_out[401];
    assign  image_1_465[111:96]    = Conv_out[400];
    assign  image_1_465[95:80]     = Conv_out[372];
    assign  image_1_465[79:64]     = Conv_out[371];
    assign  image_1_465[63:48]     = Conv_out[370];
    assign  image_1_465[47:32]     = Conv_out[342];
    assign  image_1_465[31:16]     = Conv_out[341];
    assign  image_1_465[15:0]      = Conv_out[340];

    assign  image_1_466[143:128]   = Conv_out[401];
    assign  image_1_466[127:112]   = Conv_out[400];
    assign  image_1_466[111:96]    = Conv_out[399];
    assign  image_1_466[95:80]     = Conv_out[371];
    assign  image_1_466[79:64]     = Conv_out[370];
    assign  image_1_466[63:48]     = Conv_out[369];
    assign  image_1_466[47:32]     = Conv_out[341];
    assign  image_1_466[31:16]     = Conv_out[340];
    assign  image_1_466[15:0]      = Conv_out[339];

    assign  image_1_467[143:128]   = Conv_out[400];
    assign  image_1_467[127:112]   = Conv_out[399];
    assign  image_1_467[111:96]    = Conv_out[398];
    assign  image_1_467[95:80]     = Conv_out[370];
    assign  image_1_467[79:64]     = Conv_out[369];
    assign  image_1_467[63:48]     = Conv_out[368];
    assign  image_1_467[47:32]     = Conv_out[340];
    assign  image_1_467[31:16]     = Conv_out[339];
    assign  image_1_467[15:0]      = Conv_out[338];

    assign  image_1_468[143:128]   = Conv_out[399];
    assign  image_1_468[127:112]   = Conv_out[398];
    assign  image_1_468[111:96]    = Conv_out[397];
    assign  image_1_468[95:80]     = Conv_out[369];
    assign  image_1_468[79:64]     = Conv_out[368];
    assign  image_1_468[63:48]     = Conv_out[367];
    assign  image_1_468[47:32]     = Conv_out[339];
    assign  image_1_468[31:16]     = Conv_out[338];
    assign  image_1_468[15:0]      = Conv_out[337];

    assign  image_1_469[143:128]   = Conv_out[398];
    assign  image_1_469[127:112]   = Conv_out[397];
    assign  image_1_469[111:96]    = Conv_out[396];
    assign  image_1_469[95:80]     = Conv_out[368];
    assign  image_1_469[79:64]     = Conv_out[367];
    assign  image_1_469[63:48]     = Conv_out[366];
    assign  image_1_469[47:32]     = Conv_out[338];
    assign  image_1_469[31:16]     = Conv_out[337];
    assign  image_1_469[15:0]      = Conv_out[336];

    assign  image_1_470[143:128]   = Conv_out[397];
    assign  image_1_470[127:112]   = Conv_out[396];
    assign  image_1_470[111:96]    = Conv_out[395];
    assign  image_1_470[95:80]     = Conv_out[367];
    assign  image_1_470[79:64]     = Conv_out[366];
    assign  image_1_470[63:48]     = Conv_out[365];
    assign  image_1_470[47:32]     = Conv_out[337];
    assign  image_1_470[31:16]     = Conv_out[336];
    assign  image_1_470[15:0]      = Conv_out[335];

    assign  image_1_471[143:128]   = Conv_out[396];
    assign  image_1_471[127:112]   = Conv_out[395];
    assign  image_1_471[111:96]    = Conv_out[394];
    assign  image_1_471[95:80]     = Conv_out[366];
    assign  image_1_471[79:64]     = Conv_out[365];
    assign  image_1_471[63:48]     = Conv_out[364];
    assign  image_1_471[47:32]     = Conv_out[336];
    assign  image_1_471[31:16]     = Conv_out[335];
    assign  image_1_471[15:0]      = Conv_out[334];

    assign  image_1_472[143:128]   = Conv_out[395];
    assign  image_1_472[127:112]   = Conv_out[394];
    assign  image_1_472[111:96]    = Conv_out[393];
    assign  image_1_472[95:80]     = Conv_out[365];
    assign  image_1_472[79:64]     = Conv_out[364];
    assign  image_1_472[63:48]     = Conv_out[363];
    assign  image_1_472[47:32]     = Conv_out[335];
    assign  image_1_472[31:16]     = Conv_out[334];
    assign  image_1_472[15:0]      = Conv_out[333];

    assign  image_1_473[143:128]   = Conv_out[394];
    assign  image_1_473[127:112]   = Conv_out[393];
    assign  image_1_473[111:96]    = Conv_out[392];
    assign  image_1_473[95:80]     = Conv_out[364];
    assign  image_1_473[79:64]     = Conv_out[363];
    assign  image_1_473[63:48]     = Conv_out[362];
    assign  image_1_473[47:32]     = Conv_out[334];
    assign  image_1_473[31:16]     = Conv_out[333];
    assign  image_1_473[15:0]      = Conv_out[332];

    assign  image_1_474[143:128]   = Conv_out[393];
    assign  image_1_474[127:112]   = Conv_out[392];
    assign  image_1_474[111:96]    = Conv_out[391];
    assign  image_1_474[95:80]     = Conv_out[363];
    assign  image_1_474[79:64]     = Conv_out[362];
    assign  image_1_474[63:48]     = Conv_out[361];
    assign  image_1_474[47:32]     = Conv_out[333];
    assign  image_1_474[31:16]     = Conv_out[332];
    assign  image_1_474[15:0]      = Conv_out[331];

    assign  image_1_475[143:128]   = Conv_out[392];
    assign  image_1_475[127:112]   = Conv_out[391];
    assign  image_1_475[111:96]    = Conv_out[390];
    assign  image_1_475[95:80]     = Conv_out[362];
    assign  image_1_475[79:64]     = Conv_out[361];
    assign  image_1_475[63:48]     = Conv_out[360];
    assign  image_1_475[47:32]     = Conv_out[332];
    assign  image_1_475[31:16]     = Conv_out[331];
    assign  image_1_475[15:0]      = Conv_out[330];

    assign  image_1_476[143:128]   = Conv_out[389];
    assign  image_1_476[127:112]   = Conv_out[388];
    assign  image_1_476[111:96]    = Conv_out[387];
    assign  image_1_476[95:80]     = Conv_out[359];
    assign  image_1_476[79:64]     = Conv_out[358];
    assign  image_1_476[63:48]     = Conv_out[357];
    assign  image_1_476[47:32]     = Conv_out[329];
    assign  image_1_476[31:16]     = Conv_out[328];
    assign  image_1_476[15:0]      = Conv_out[327];

    assign  image_1_477[143:128]   = Conv_out[388];
    assign  image_1_477[127:112]   = Conv_out[387];
    assign  image_1_477[111:96]    = Conv_out[386];
    assign  image_1_477[95:80]     = Conv_out[358];
    assign  image_1_477[79:64]     = Conv_out[357];
    assign  image_1_477[63:48]     = Conv_out[356];
    assign  image_1_477[47:32]     = Conv_out[328];
    assign  image_1_477[31:16]     = Conv_out[327];
    assign  image_1_477[15:0]      = Conv_out[326];

    assign  image_1_478[143:128]   = Conv_out[387];
    assign  image_1_478[127:112]   = Conv_out[386];
    assign  image_1_478[111:96]    = Conv_out[385];
    assign  image_1_478[95:80]     = Conv_out[357];
    assign  image_1_478[79:64]     = Conv_out[356];
    assign  image_1_478[63:48]     = Conv_out[355];
    assign  image_1_478[47:32]     = Conv_out[327];
    assign  image_1_478[31:16]     = Conv_out[326];
    assign  image_1_478[15:0]      = Conv_out[325];

    assign  image_1_479[143:128]   = Conv_out[386];
    assign  image_1_479[127:112]   = Conv_out[385];
    assign  image_1_479[111:96]    = Conv_out[384];
    assign  image_1_479[95:80]     = Conv_out[356];
    assign  image_1_479[79:64]     = Conv_out[355];
    assign  image_1_479[63:48]     = Conv_out[354];
    assign  image_1_479[47:32]     = Conv_out[326];
    assign  image_1_479[31:16]     = Conv_out[325];
    assign  image_1_479[15:0]      = Conv_out[324];

    assign  image_1_480[143:128]   = Conv_out[385];
    assign  image_1_480[127:112]   = Conv_out[384];
    assign  image_1_480[111:96]    = Conv_out[383];
    assign  image_1_480[95:80]     = Conv_out[355];
    assign  image_1_480[79:64]     = Conv_out[354];
    assign  image_1_480[63:48]     = Conv_out[353];
    assign  image_1_480[47:32]     = Conv_out[325];
    assign  image_1_480[31:16]     = Conv_out[324];
    assign  image_1_480[15:0]      = Conv_out[323];

    assign  image_1_481[143:128]   = Conv_out[384];
    assign  image_1_481[127:112]   = Conv_out[383];
    assign  image_1_481[111:96]    = Conv_out[382];
    assign  image_1_481[95:80]     = Conv_out[354];
    assign  image_1_481[79:64]     = Conv_out[353];
    assign  image_1_481[63:48]     = Conv_out[352];
    assign  image_1_481[47:32]     = Conv_out[324];
    assign  image_1_481[31:16]     = Conv_out[323];
    assign  image_1_481[15:0]      = Conv_out[322];

    assign  image_1_482[143:128]   = Conv_out[383];
    assign  image_1_482[127:112]   = Conv_out[382];
    assign  image_1_482[111:96]    = Conv_out[381];
    assign  image_1_482[95:80]     = Conv_out[353];
    assign  image_1_482[79:64]     = Conv_out[352];
    assign  image_1_482[63:48]     = Conv_out[351];
    assign  image_1_482[47:32]     = Conv_out[323];
    assign  image_1_482[31:16]     = Conv_out[322];
    assign  image_1_482[15:0]      = Conv_out[321];

    assign  image_1_483[143:128]   = Conv_out[382];
    assign  image_1_483[127:112]   = Conv_out[381];
    assign  image_1_483[111:96]    = Conv_out[380];
    assign  image_1_483[95:80]     = Conv_out[352];
    assign  image_1_483[79:64]     = Conv_out[351];
    assign  image_1_483[63:48]     = Conv_out[350];
    assign  image_1_483[47:32]     = Conv_out[322];
    assign  image_1_483[31:16]     = Conv_out[321];
    assign  image_1_483[15:0]      = Conv_out[320];

    assign  image_1_484[143:128]   = Conv_out[381];
    assign  image_1_484[127:112]   = Conv_out[380];
    assign  image_1_484[111:96]    = Conv_out[379];
    assign  image_1_484[95:80]     = Conv_out[351];
    assign  image_1_484[79:64]     = Conv_out[350];
    assign  image_1_484[63:48]     = Conv_out[349];
    assign  image_1_484[47:32]     = Conv_out[321];
    assign  image_1_484[31:16]     = Conv_out[320];
    assign  image_1_484[15:0]      = Conv_out[319];

    assign  image_1_485[143:128]   = Conv_out[380];
    assign  image_1_485[127:112]   = Conv_out[379];
    assign  image_1_485[111:96]    = Conv_out[378];
    assign  image_1_485[95:80]     = Conv_out[350];
    assign  image_1_485[79:64]     = Conv_out[349];
    assign  image_1_485[63:48]     = Conv_out[348];
    assign  image_1_485[47:32]     = Conv_out[320];
    assign  image_1_485[31:16]     = Conv_out[319];
    assign  image_1_485[15:0]      = Conv_out[318];

    assign  image_1_486[143:128]   = Conv_out[379];
    assign  image_1_486[127:112]   = Conv_out[378];
    assign  image_1_486[111:96]    = Conv_out[377];
    assign  image_1_486[95:80]     = Conv_out[349];
    assign  image_1_486[79:64]     = Conv_out[348];
    assign  image_1_486[63:48]     = Conv_out[347];
    assign  image_1_486[47:32]     = Conv_out[319];
    assign  image_1_486[31:16]     = Conv_out[318];
    assign  image_1_486[15:0]      = Conv_out[317];

    assign  image_1_487[143:128]   = Conv_out[378];
    assign  image_1_487[127:112]   = Conv_out[377];
    assign  image_1_487[111:96]    = Conv_out[376];
    assign  image_1_487[95:80]     = Conv_out[348];
    assign  image_1_487[79:64]     = Conv_out[347];
    assign  image_1_487[63:48]     = Conv_out[346];
    assign  image_1_487[47:32]     = Conv_out[318];
    assign  image_1_487[31:16]     = Conv_out[317];
    assign  image_1_487[15:0]      = Conv_out[316];

    assign  image_1_488[143:128]   = Conv_out[377];
    assign  image_1_488[127:112]   = Conv_out[376];
    assign  image_1_488[111:96]    = Conv_out[375];
    assign  image_1_488[95:80]     = Conv_out[347];
    assign  image_1_488[79:64]     = Conv_out[346];
    assign  image_1_488[63:48]     = Conv_out[345];
    assign  image_1_488[47:32]     = Conv_out[317];
    assign  image_1_488[31:16]     = Conv_out[316];
    assign  image_1_488[15:0]      = Conv_out[315];

    assign  image_1_489[143:128]   = Conv_out[376];
    assign  image_1_489[127:112]   = Conv_out[375];
    assign  image_1_489[111:96]    = Conv_out[374];
    assign  image_1_489[95:80]     = Conv_out[346];
    assign  image_1_489[79:64]     = Conv_out[345];
    assign  image_1_489[63:48]     = Conv_out[344];
    assign  image_1_489[47:32]     = Conv_out[316];
    assign  image_1_489[31:16]     = Conv_out[315];
    assign  image_1_489[15:0]      = Conv_out[314];

    assign  image_1_490[143:128]   = Conv_out[375];
    assign  image_1_490[127:112]   = Conv_out[374];
    assign  image_1_490[111:96]    = Conv_out[373];
    assign  image_1_490[95:80]     = Conv_out[345];
    assign  image_1_490[79:64]     = Conv_out[344];
    assign  image_1_490[63:48]     = Conv_out[343];
    assign  image_1_490[47:32]     = Conv_out[315];
    assign  image_1_490[31:16]     = Conv_out[314];
    assign  image_1_490[15:0]      = Conv_out[313];

    assign  image_1_491[143:128]   = Conv_out[374];
    assign  image_1_491[127:112]   = Conv_out[373];
    assign  image_1_491[111:96]    = Conv_out[372];
    assign  image_1_491[95:80]     = Conv_out[344];
    assign  image_1_491[79:64]     = Conv_out[343];
    assign  image_1_491[63:48]     = Conv_out[342];
    assign  image_1_491[47:32]     = Conv_out[314];
    assign  image_1_491[31:16]     = Conv_out[313];
    assign  image_1_491[15:0]      = Conv_out[312];

    assign  image_1_492[143:128]   = Conv_out[373];
    assign  image_1_492[127:112]   = Conv_out[372];
    assign  image_1_492[111:96]    = Conv_out[371];
    assign  image_1_492[95:80]     = Conv_out[343];
    assign  image_1_492[79:64]     = Conv_out[342];
    assign  image_1_492[63:48]     = Conv_out[341];
    assign  image_1_492[47:32]     = Conv_out[313];
    assign  image_1_492[31:16]     = Conv_out[312];
    assign  image_1_492[15:0]      = Conv_out[311];

    assign  image_1_493[143:128]   = Conv_out[372];
    assign  image_1_493[127:112]   = Conv_out[371];
    assign  image_1_493[111:96]    = Conv_out[370];
    assign  image_1_493[95:80]     = Conv_out[342];
    assign  image_1_493[79:64]     = Conv_out[341];
    assign  image_1_493[63:48]     = Conv_out[340];
    assign  image_1_493[47:32]     = Conv_out[312];
    assign  image_1_493[31:16]     = Conv_out[311];
    assign  image_1_493[15:0]      = Conv_out[310];

    assign  image_1_494[143:128]   = Conv_out[371];
    assign  image_1_494[127:112]   = Conv_out[370];
    assign  image_1_494[111:96]    = Conv_out[369];
    assign  image_1_494[95:80]     = Conv_out[341];
    assign  image_1_494[79:64]     = Conv_out[340];
    assign  image_1_494[63:48]     = Conv_out[339];
    assign  image_1_494[47:32]     = Conv_out[311];
    assign  image_1_494[31:16]     = Conv_out[310];
    assign  image_1_494[15:0]      = Conv_out[309];

    assign  image_1_495[143:128]   = Conv_out[370];
    assign  image_1_495[127:112]   = Conv_out[369];
    assign  image_1_495[111:96]    = Conv_out[368];
    assign  image_1_495[95:80]     = Conv_out[340];
    assign  image_1_495[79:64]     = Conv_out[339];
    assign  image_1_495[63:48]     = Conv_out[338];
    assign  image_1_495[47:32]     = Conv_out[310];
    assign  image_1_495[31:16]     = Conv_out[309];
    assign  image_1_495[15:0]      = Conv_out[308];

    assign  image_1_496[143:128]   = Conv_out[369];
    assign  image_1_496[127:112]   = Conv_out[368];
    assign  image_1_496[111:96]    = Conv_out[367];
    assign  image_1_496[95:80]     = Conv_out[339];
    assign  image_1_496[79:64]     = Conv_out[338];
    assign  image_1_496[63:48]     = Conv_out[337];
    assign  image_1_496[47:32]     = Conv_out[309];
    assign  image_1_496[31:16]     = Conv_out[308];
    assign  image_1_496[15:0]      = Conv_out[307];

    assign  image_1_497[143:128]   = Conv_out[368];
    assign  image_1_497[127:112]   = Conv_out[367];
    assign  image_1_497[111:96]    = Conv_out[366];
    assign  image_1_497[95:80]     = Conv_out[338];
    assign  image_1_497[79:64]     = Conv_out[337];
    assign  image_1_497[63:48]     = Conv_out[336];
    assign  image_1_497[47:32]     = Conv_out[308];
    assign  image_1_497[31:16]     = Conv_out[307];
    assign  image_1_497[15:0]      = Conv_out[306];

    assign  image_1_498[143:128]   = Conv_out[367];
    assign  image_1_498[127:112]   = Conv_out[366];
    assign  image_1_498[111:96]    = Conv_out[365];
    assign  image_1_498[95:80]     = Conv_out[337];
    assign  image_1_498[79:64]     = Conv_out[336];
    assign  image_1_498[63:48]     = Conv_out[335];
    assign  image_1_498[47:32]     = Conv_out[307];
    assign  image_1_498[31:16]     = Conv_out[306];
    assign  image_1_498[15:0]      = Conv_out[305];

    assign  image_1_499[143:128]   = Conv_out[366];
    assign  image_1_499[127:112]   = Conv_out[365];
    assign  image_1_499[111:96]    = Conv_out[364];
    assign  image_1_499[95:80]     = Conv_out[336];
    assign  image_1_499[79:64]     = Conv_out[335];
    assign  image_1_499[63:48]     = Conv_out[334];
    assign  image_1_499[47:32]     = Conv_out[306];
    assign  image_1_499[31:16]     = Conv_out[305];
    assign  image_1_499[15:0]      = Conv_out[304];

    assign  image_1_500[143:128]   = Conv_out[365];
    assign  image_1_500[127:112]   = Conv_out[364];
    assign  image_1_500[111:96]    = Conv_out[363];
    assign  image_1_500[95:80]     = Conv_out[335];
    assign  image_1_500[79:64]     = Conv_out[334];
    assign  image_1_500[63:48]     = Conv_out[333];
    assign  image_1_500[47:32]     = Conv_out[305];
    assign  image_1_500[31:16]     = Conv_out[304];
    assign  image_1_500[15:0]      = Conv_out[303];

    assign  image_1_501[143:128]   = Conv_out[364];
    assign  image_1_501[127:112]   = Conv_out[363];
    assign  image_1_501[111:96]    = Conv_out[362];
    assign  image_1_501[95:80]     = Conv_out[334];
    assign  image_1_501[79:64]     = Conv_out[333];
    assign  image_1_501[63:48]     = Conv_out[332];
    assign  image_1_501[47:32]     = Conv_out[304];
    assign  image_1_501[31:16]     = Conv_out[303];
    assign  image_1_501[15:0]      = Conv_out[302];

    assign  image_1_502[143:128]   = Conv_out[363];
    assign  image_1_502[127:112]   = Conv_out[362];
    assign  image_1_502[111:96]    = Conv_out[361];
    assign  image_1_502[95:80]     = Conv_out[333];
    assign  image_1_502[79:64]     = Conv_out[332];
    assign  image_1_502[63:48]     = Conv_out[331];
    assign  image_1_502[47:32]     = Conv_out[303];
    assign  image_1_502[31:16]     = Conv_out[302];
    assign  image_1_502[15:0]      = Conv_out[301];

    assign  image_1_503[143:128]   = Conv_out[362];
    assign  image_1_503[127:112]   = Conv_out[361];
    assign  image_1_503[111:96]    = Conv_out[360];
    assign  image_1_503[95:80]     = Conv_out[332];
    assign  image_1_503[79:64]     = Conv_out[331];
    assign  image_1_503[63:48]     = Conv_out[330];
    assign  image_1_503[47:32]     = Conv_out[302];
    assign  image_1_503[31:16]     = Conv_out[301];
    assign  image_1_503[15:0]      = Conv_out[300];

    assign  image_1_504[143:128]   = Conv_out[359];
    assign  image_1_504[127:112]   = Conv_out[358];
    assign  image_1_504[111:96]    = Conv_out[357];
    assign  image_1_504[95:80]     = Conv_out[329];
    assign  image_1_504[79:64]     = Conv_out[328];
    assign  image_1_504[63:48]     = Conv_out[327];
    assign  image_1_504[47:32]     = Conv_out[299];
    assign  image_1_504[31:16]     = Conv_out[298];
    assign  image_1_504[15:0]      = Conv_out[297];

    assign  image_1_505[143:128]   = Conv_out[358];
    assign  image_1_505[127:112]   = Conv_out[357];
    assign  image_1_505[111:96]    = Conv_out[356];
    assign  image_1_505[95:80]     = Conv_out[328];
    assign  image_1_505[79:64]     = Conv_out[327];
    assign  image_1_505[63:48]     = Conv_out[326];
    assign  image_1_505[47:32]     = Conv_out[298];
    assign  image_1_505[31:16]     = Conv_out[297];
    assign  image_1_505[15:0]      = Conv_out[296];

    assign  image_1_506[143:128]   = Conv_out[357];
    assign  image_1_506[127:112]   = Conv_out[356];
    assign  image_1_506[111:96]    = Conv_out[355];
    assign  image_1_506[95:80]     = Conv_out[327];
    assign  image_1_506[79:64]     = Conv_out[326];
    assign  image_1_506[63:48]     = Conv_out[325];
    assign  image_1_506[47:32]     = Conv_out[297];
    assign  image_1_506[31:16]     = Conv_out[296];
    assign  image_1_506[15:0]      = Conv_out[295];

    assign  image_1_507[143:128]   = Conv_out[356];
    assign  image_1_507[127:112]   = Conv_out[355];
    assign  image_1_507[111:96]    = Conv_out[354];
    assign  image_1_507[95:80]     = Conv_out[326];
    assign  image_1_507[79:64]     = Conv_out[325];
    assign  image_1_507[63:48]     = Conv_out[324];
    assign  image_1_507[47:32]     = Conv_out[296];
    assign  image_1_507[31:16]     = Conv_out[295];
    assign  image_1_507[15:0]      = Conv_out[294];

    assign  image_1_508[143:128]   = Conv_out[355];
    assign  image_1_508[127:112]   = Conv_out[354];
    assign  image_1_508[111:96]    = Conv_out[353];
    assign  image_1_508[95:80]     = Conv_out[325];
    assign  image_1_508[79:64]     = Conv_out[324];
    assign  image_1_508[63:48]     = Conv_out[323];
    assign  image_1_508[47:32]     = Conv_out[295];
    assign  image_1_508[31:16]     = Conv_out[294];
    assign  image_1_508[15:0]      = Conv_out[293];

    assign  image_1_509[143:128]   = Conv_out[354];
    assign  image_1_509[127:112]   = Conv_out[353];
    assign  image_1_509[111:96]    = Conv_out[352];
    assign  image_1_509[95:80]     = Conv_out[324];
    assign  image_1_509[79:64]     = Conv_out[323];
    assign  image_1_509[63:48]     = Conv_out[322];
    assign  image_1_509[47:32]     = Conv_out[294];
    assign  image_1_509[31:16]     = Conv_out[293];
    assign  image_1_509[15:0]      = Conv_out[292];

    assign  image_1_510[143:128]   = Conv_out[353];
    assign  image_1_510[127:112]   = Conv_out[352];
    assign  image_1_510[111:96]    = Conv_out[351];
    assign  image_1_510[95:80]     = Conv_out[323];
    assign  image_1_510[79:64]     = Conv_out[322];
    assign  image_1_510[63:48]     = Conv_out[321];
    assign  image_1_510[47:32]     = Conv_out[293];
    assign  image_1_510[31:16]     = Conv_out[292];
    assign  image_1_510[15:0]      = Conv_out[291];

    assign  image_1_511[143:128]   = Conv_out[352];
    assign  image_1_511[127:112]   = Conv_out[351];
    assign  image_1_511[111:96]    = Conv_out[350];
    assign  image_1_511[95:80]     = Conv_out[322];
    assign  image_1_511[79:64]     = Conv_out[321];
    assign  image_1_511[63:48]     = Conv_out[320];
    assign  image_1_511[47:32]     = Conv_out[292];
    assign  image_1_511[31:16]     = Conv_out[291];
    assign  image_1_511[15:0]      = Conv_out[290];

    assign  image_1_512[143:128]   = Conv_out[351];
    assign  image_1_512[127:112]   = Conv_out[350];
    assign  image_1_512[111:96]    = Conv_out[349];
    assign  image_1_512[95:80]     = Conv_out[321];
    assign  image_1_512[79:64]     = Conv_out[320];
    assign  image_1_512[63:48]     = Conv_out[319];
    assign  image_1_512[47:32]     = Conv_out[291];
    assign  image_1_512[31:16]     = Conv_out[290];
    assign  image_1_512[15:0]      = Conv_out[289];

    assign  image_1_513[143:128]   = Conv_out[350];
    assign  image_1_513[127:112]   = Conv_out[349];
    assign  image_1_513[111:96]    = Conv_out[348];
    assign  image_1_513[95:80]     = Conv_out[320];
    assign  image_1_513[79:64]     = Conv_out[319];
    assign  image_1_513[63:48]     = Conv_out[318];
    assign  image_1_513[47:32]     = Conv_out[290];
    assign  image_1_513[31:16]     = Conv_out[289];
    assign  image_1_513[15:0]      = Conv_out[288];

    assign  image_1_514[143:128]   = Conv_out[349];
    assign  image_1_514[127:112]   = Conv_out[348];
    assign  image_1_514[111:96]    = Conv_out[347];
    assign  image_1_514[95:80]     = Conv_out[319];
    assign  image_1_514[79:64]     = Conv_out[318];
    assign  image_1_514[63:48]     = Conv_out[317];
    assign  image_1_514[47:32]     = Conv_out[289];
    assign  image_1_514[31:16]     = Conv_out[288];
    assign  image_1_514[15:0]      = Conv_out[287];

    assign  image_1_515[143:128]   = Conv_out[348];
    assign  image_1_515[127:112]   = Conv_out[347];
    assign  image_1_515[111:96]    = Conv_out[346];
    assign  image_1_515[95:80]     = Conv_out[318];
    assign  image_1_515[79:64]     = Conv_out[317];
    assign  image_1_515[63:48]     = Conv_out[316];
    assign  image_1_515[47:32]     = Conv_out[288];
    assign  image_1_515[31:16]     = Conv_out[287];
    assign  image_1_515[15:0]      = Conv_out[286];

    assign  image_1_516[143:128]   = Conv_out[347];
    assign  image_1_516[127:112]   = Conv_out[346];
    assign  image_1_516[111:96]    = Conv_out[345];
    assign  image_1_516[95:80]     = Conv_out[317];
    assign  image_1_516[79:64]     = Conv_out[316];
    assign  image_1_516[63:48]     = Conv_out[315];
    assign  image_1_516[47:32]     = Conv_out[287];
    assign  image_1_516[31:16]     = Conv_out[286];
    assign  image_1_516[15:0]      = Conv_out[285];

    assign  image_1_517[143:128]   = Conv_out[346];
    assign  image_1_517[127:112]   = Conv_out[345];
    assign  image_1_517[111:96]    = Conv_out[344];
    assign  image_1_517[95:80]     = Conv_out[316];
    assign  image_1_517[79:64]     = Conv_out[315];
    assign  image_1_517[63:48]     = Conv_out[314];
    assign  image_1_517[47:32]     = Conv_out[286];
    assign  image_1_517[31:16]     = Conv_out[285];
    assign  image_1_517[15:0]      = Conv_out[284];

    assign  image_1_518[143:128]   = Conv_out[345];
    assign  image_1_518[127:112]   = Conv_out[344];
    assign  image_1_518[111:96]    = Conv_out[343];
    assign  image_1_518[95:80]     = Conv_out[315];
    assign  image_1_518[79:64]     = Conv_out[314];
    assign  image_1_518[63:48]     = Conv_out[313];
    assign  image_1_518[47:32]     = Conv_out[285];
    assign  image_1_518[31:16]     = Conv_out[284];
    assign  image_1_518[15:0]      = Conv_out[283];

    assign  image_1_519[143:128]   = Conv_out[344];
    assign  image_1_519[127:112]   = Conv_out[343];
    assign  image_1_519[111:96]    = Conv_out[342];
    assign  image_1_519[95:80]     = Conv_out[314];
    assign  image_1_519[79:64]     = Conv_out[313];
    assign  image_1_519[63:48]     = Conv_out[312];
    assign  image_1_519[47:32]     = Conv_out[284];
    assign  image_1_519[31:16]     = Conv_out[283];
    assign  image_1_519[15:0]      = Conv_out[282];

    assign  image_1_520[143:128]   = Conv_out[343];
    assign  image_1_520[127:112]   = Conv_out[342];
    assign  image_1_520[111:96]    = Conv_out[341];
    assign  image_1_520[95:80]     = Conv_out[313];
    assign  image_1_520[79:64]     = Conv_out[312];
    assign  image_1_520[63:48]     = Conv_out[311];
    assign  image_1_520[47:32]     = Conv_out[283];
    assign  image_1_520[31:16]     = Conv_out[282];
    assign  image_1_520[15:0]      = Conv_out[281];

    assign  image_1_521[143:128]   = Conv_out[342];
    assign  image_1_521[127:112]   = Conv_out[341];
    assign  image_1_521[111:96]    = Conv_out[340];
    assign  image_1_521[95:80]     = Conv_out[312];
    assign  image_1_521[79:64]     = Conv_out[311];
    assign  image_1_521[63:48]     = Conv_out[310];
    assign  image_1_521[47:32]     = Conv_out[282];
    assign  image_1_521[31:16]     = Conv_out[281];
    assign  image_1_521[15:0]      = Conv_out[280];

    assign  image_1_522[143:128]   = Conv_out[341];
    assign  image_1_522[127:112]   = Conv_out[340];
    assign  image_1_522[111:96]    = Conv_out[339];
    assign  image_1_522[95:80]     = Conv_out[311];
    assign  image_1_522[79:64]     = Conv_out[310];
    assign  image_1_522[63:48]     = Conv_out[309];
    assign  image_1_522[47:32]     = Conv_out[281];
    assign  image_1_522[31:16]     = Conv_out[280];
    assign  image_1_522[15:0]      = Conv_out[279];

    assign  image_1_523[143:128]   = Conv_out[340];
    assign  image_1_523[127:112]   = Conv_out[339];
    assign  image_1_523[111:96]    = Conv_out[338];
    assign  image_1_523[95:80]     = Conv_out[310];
    assign  image_1_523[79:64]     = Conv_out[309];
    assign  image_1_523[63:48]     = Conv_out[308];
    assign  image_1_523[47:32]     = Conv_out[280];
    assign  image_1_523[31:16]     = Conv_out[279];
    assign  image_1_523[15:0]      = Conv_out[278];

    assign  image_1_524[143:128]   = Conv_out[339];
    assign  image_1_524[127:112]   = Conv_out[338];
    assign  image_1_524[111:96]    = Conv_out[337];
    assign  image_1_524[95:80]     = Conv_out[309];
    assign  image_1_524[79:64]     = Conv_out[308];
    assign  image_1_524[63:48]     = Conv_out[307];
    assign  image_1_524[47:32]     = Conv_out[279];
    assign  image_1_524[31:16]     = Conv_out[278];
    assign  image_1_524[15:0]      = Conv_out[277];

    assign  image_1_525[143:128]   = Conv_out[338];
    assign  image_1_525[127:112]   = Conv_out[337];
    assign  image_1_525[111:96]    = Conv_out[336];
    assign  image_1_525[95:80]     = Conv_out[308];
    assign  image_1_525[79:64]     = Conv_out[307];
    assign  image_1_525[63:48]     = Conv_out[306];
    assign  image_1_525[47:32]     = Conv_out[278];
    assign  image_1_525[31:16]     = Conv_out[277];
    assign  image_1_525[15:0]      = Conv_out[276];

    assign  image_1_526[143:128]   = Conv_out[337];
    assign  image_1_526[127:112]   = Conv_out[336];
    assign  image_1_526[111:96]    = Conv_out[335];
    assign  image_1_526[95:80]     = Conv_out[307];
    assign  image_1_526[79:64]     = Conv_out[306];
    assign  image_1_526[63:48]     = Conv_out[305];
    assign  image_1_526[47:32]     = Conv_out[277];
    assign  image_1_526[31:16]     = Conv_out[276];
    assign  image_1_526[15:0]      = Conv_out[275];

    assign  image_1_527[143:128]   = Conv_out[336];
    assign  image_1_527[127:112]   = Conv_out[335];
    assign  image_1_527[111:96]    = Conv_out[334];
    assign  image_1_527[95:80]     = Conv_out[306];
    assign  image_1_527[79:64]     = Conv_out[305];
    assign  image_1_527[63:48]     = Conv_out[304];
    assign  image_1_527[47:32]     = Conv_out[276];
    assign  image_1_527[31:16]     = Conv_out[275];
    assign  image_1_527[15:0]      = Conv_out[274];

    assign  image_1_528[143:128]   = Conv_out[335];
    assign  image_1_528[127:112]   = Conv_out[334];
    assign  image_1_528[111:96]    = Conv_out[333];
    assign  image_1_528[95:80]     = Conv_out[305];
    assign  image_1_528[79:64]     = Conv_out[304];
    assign  image_1_528[63:48]     = Conv_out[303];
    assign  image_1_528[47:32]     = Conv_out[275];
    assign  image_1_528[31:16]     = Conv_out[274];
    assign  image_1_528[15:0]      = Conv_out[273];

    assign  image_1_529[143:128]   = Conv_out[334];
    assign  image_1_529[127:112]   = Conv_out[333];
    assign  image_1_529[111:96]    = Conv_out[332];
    assign  image_1_529[95:80]     = Conv_out[304];
    assign  image_1_529[79:64]     = Conv_out[303];
    assign  image_1_529[63:48]     = Conv_out[302];
    assign  image_1_529[47:32]     = Conv_out[274];
    assign  image_1_529[31:16]     = Conv_out[273];
    assign  image_1_529[15:0]      = Conv_out[272];

    assign  image_1_530[143:128]   = Conv_out[333];
    assign  image_1_530[127:112]   = Conv_out[332];
    assign  image_1_530[111:96]    = Conv_out[331];
    assign  image_1_530[95:80]     = Conv_out[303];
    assign  image_1_530[79:64]     = Conv_out[302];
    assign  image_1_530[63:48]     = Conv_out[301];
    assign  image_1_530[47:32]     = Conv_out[273];
    assign  image_1_530[31:16]     = Conv_out[272];
    assign  image_1_530[15:0]      = Conv_out[271];

    assign  image_1_531[143:128]   = Conv_out[332];
    assign  image_1_531[127:112]   = Conv_out[331];
    assign  image_1_531[111:96]    = Conv_out[330];
    assign  image_1_531[95:80]     = Conv_out[302];
    assign  image_1_531[79:64]     = Conv_out[301];
    assign  image_1_531[63:48]     = Conv_out[300];
    assign  image_1_531[47:32]     = Conv_out[272];
    assign  image_1_531[31:16]     = Conv_out[271];
    assign  image_1_531[15:0]      = Conv_out[270];

    assign  image_1_532[143:128]   = Conv_out[329];
    assign  image_1_532[127:112]   = Conv_out[328];
    assign  image_1_532[111:96]    = Conv_out[327];
    assign  image_1_532[95:80]     = Conv_out[299];
    assign  image_1_532[79:64]     = Conv_out[298];
    assign  image_1_532[63:48]     = Conv_out[297];
    assign  image_1_532[47:32]     = Conv_out[269];
    assign  image_1_532[31:16]     = Conv_out[268];
    assign  image_1_532[15:0]      = Conv_out[267];

    assign  image_1_533[143:128]   = Conv_out[328];
    assign  image_1_533[127:112]   = Conv_out[327];
    assign  image_1_533[111:96]    = Conv_out[326];
    assign  image_1_533[95:80]     = Conv_out[298];
    assign  image_1_533[79:64]     = Conv_out[297];
    assign  image_1_533[63:48]     = Conv_out[296];
    assign  image_1_533[47:32]     = Conv_out[268];
    assign  image_1_533[31:16]     = Conv_out[267];
    assign  image_1_533[15:0]      = Conv_out[266];

    assign  image_1_534[143:128]   = Conv_out[327];
    assign  image_1_534[127:112]   = Conv_out[326];
    assign  image_1_534[111:96]    = Conv_out[325];
    assign  image_1_534[95:80]     = Conv_out[297];
    assign  image_1_534[79:64]     = Conv_out[296];
    assign  image_1_534[63:48]     = Conv_out[295];
    assign  image_1_534[47:32]     = Conv_out[267];
    assign  image_1_534[31:16]     = Conv_out[266];
    assign  image_1_534[15:0]      = Conv_out[265];

    assign  image_1_535[143:128]   = Conv_out[326];
    assign  image_1_535[127:112]   = Conv_out[325];
    assign  image_1_535[111:96]    = Conv_out[324];
    assign  image_1_535[95:80]     = Conv_out[296];
    assign  image_1_535[79:64]     = Conv_out[295];
    assign  image_1_535[63:48]     = Conv_out[294];
    assign  image_1_535[47:32]     = Conv_out[266];
    assign  image_1_535[31:16]     = Conv_out[265];
    assign  image_1_535[15:0]      = Conv_out[264];

    assign  image_1_536[143:128]   = Conv_out[325];
    assign  image_1_536[127:112]   = Conv_out[324];
    assign  image_1_536[111:96]    = Conv_out[323];
    assign  image_1_536[95:80]     = Conv_out[295];
    assign  image_1_536[79:64]     = Conv_out[294];
    assign  image_1_536[63:48]     = Conv_out[293];
    assign  image_1_536[47:32]     = Conv_out[265];
    assign  image_1_536[31:16]     = Conv_out[264];
    assign  image_1_536[15:0]      = Conv_out[263];

    assign  image_1_537[143:128]   = Conv_out[324];
    assign  image_1_537[127:112]   = Conv_out[323];
    assign  image_1_537[111:96]    = Conv_out[322];
    assign  image_1_537[95:80]     = Conv_out[294];
    assign  image_1_537[79:64]     = Conv_out[293];
    assign  image_1_537[63:48]     = Conv_out[292];
    assign  image_1_537[47:32]     = Conv_out[264];
    assign  image_1_537[31:16]     = Conv_out[263];
    assign  image_1_537[15:0]      = Conv_out[262];

    assign  image_1_538[143:128]   = Conv_out[323];
    assign  image_1_538[127:112]   = Conv_out[322];
    assign  image_1_538[111:96]    = Conv_out[321];
    assign  image_1_538[95:80]     = Conv_out[293];
    assign  image_1_538[79:64]     = Conv_out[292];
    assign  image_1_538[63:48]     = Conv_out[291];
    assign  image_1_538[47:32]     = Conv_out[263];
    assign  image_1_538[31:16]     = Conv_out[262];
    assign  image_1_538[15:0]      = Conv_out[261];

    assign  image_1_539[143:128]   = Conv_out[322];
    assign  image_1_539[127:112]   = Conv_out[321];
    assign  image_1_539[111:96]    = Conv_out[320];
    assign  image_1_539[95:80]     = Conv_out[292];
    assign  image_1_539[79:64]     = Conv_out[291];
    assign  image_1_539[63:48]     = Conv_out[290];
    assign  image_1_539[47:32]     = Conv_out[262];
    assign  image_1_539[31:16]     = Conv_out[261];
    assign  image_1_539[15:0]      = Conv_out[260];

    assign  image_1_540[143:128]   = Conv_out[321];
    assign  image_1_540[127:112]   = Conv_out[320];
    assign  image_1_540[111:96]    = Conv_out[319];
    assign  image_1_540[95:80]     = Conv_out[291];
    assign  image_1_540[79:64]     = Conv_out[290];
    assign  image_1_540[63:48]     = Conv_out[289];
    assign  image_1_540[47:32]     = Conv_out[261];
    assign  image_1_540[31:16]     = Conv_out[260];
    assign  image_1_540[15:0]      = Conv_out[259];

    assign  image_1_541[143:128]   = Conv_out[320];
    assign  image_1_541[127:112]   = Conv_out[319];
    assign  image_1_541[111:96]    = Conv_out[318];
    assign  image_1_541[95:80]     = Conv_out[290];
    assign  image_1_541[79:64]     = Conv_out[289];
    assign  image_1_541[63:48]     = Conv_out[288];
    assign  image_1_541[47:32]     = Conv_out[260];
    assign  image_1_541[31:16]     = Conv_out[259];
    assign  image_1_541[15:0]      = Conv_out[258];

    assign  image_1_542[143:128]   = Conv_out[319];
    assign  image_1_542[127:112]   = Conv_out[318];
    assign  image_1_542[111:96]    = Conv_out[317];
    assign  image_1_542[95:80]     = Conv_out[289];
    assign  image_1_542[79:64]     = Conv_out[288];
    assign  image_1_542[63:48]     = Conv_out[287];
    assign  image_1_542[47:32]     = Conv_out[259];
    assign  image_1_542[31:16]     = Conv_out[258];
    assign  image_1_542[15:0]      = Conv_out[257];

    assign  image_1_543[143:128]   = Conv_out[318];
    assign  image_1_543[127:112]   = Conv_out[317];
    assign  image_1_543[111:96]    = Conv_out[316];
    assign  image_1_543[95:80]     = Conv_out[288];
    assign  image_1_543[79:64]     = Conv_out[287];
    assign  image_1_543[63:48]     = Conv_out[286];
    assign  image_1_543[47:32]     = Conv_out[258];
    assign  image_1_543[31:16]     = Conv_out[257];
    assign  image_1_543[15:0]      = Conv_out[256];

    assign  image_1_544[143:128]   = Conv_out[317];
    assign  image_1_544[127:112]   = Conv_out[316];
    assign  image_1_544[111:96]    = Conv_out[315];
    assign  image_1_544[95:80]     = Conv_out[287];
    assign  image_1_544[79:64]     = Conv_out[286];
    assign  image_1_544[63:48]     = Conv_out[285];
    assign  image_1_544[47:32]     = Conv_out[257];
    assign  image_1_544[31:16]     = Conv_out[256];
    assign  image_1_544[15:0]      = Conv_out[255];

    assign  image_1_545[143:128]   = Conv_out[316];
    assign  image_1_545[127:112]   = Conv_out[315];
    assign  image_1_545[111:96]    = Conv_out[314];
    assign  image_1_545[95:80]     = Conv_out[286];
    assign  image_1_545[79:64]     = Conv_out[285];
    assign  image_1_545[63:48]     = Conv_out[284];
    assign  image_1_545[47:32]     = Conv_out[256];
    assign  image_1_545[31:16]     = Conv_out[255];
    assign  image_1_545[15:0]      = Conv_out[254];

    assign  image_1_546[143:128]   = Conv_out[315];
    assign  image_1_546[127:112]   = Conv_out[314];
    assign  image_1_546[111:96]    = Conv_out[313];
    assign  image_1_546[95:80]     = Conv_out[285];
    assign  image_1_546[79:64]     = Conv_out[284];
    assign  image_1_546[63:48]     = Conv_out[283];
    assign  image_1_546[47:32]     = Conv_out[255];
    assign  image_1_546[31:16]     = Conv_out[254];
    assign  image_1_546[15:0]      = Conv_out[253];

    assign  image_1_547[143:128]   = Conv_out[314];
    assign  image_1_547[127:112]   = Conv_out[313];
    assign  image_1_547[111:96]    = Conv_out[312];
    assign  image_1_547[95:80]     = Conv_out[284];
    assign  image_1_547[79:64]     = Conv_out[283];
    assign  image_1_547[63:48]     = Conv_out[282];
    assign  image_1_547[47:32]     = Conv_out[254];
    assign  image_1_547[31:16]     = Conv_out[253];
    assign  image_1_547[15:0]      = Conv_out[252];

    assign  image_1_548[143:128]   = Conv_out[313];
    assign  image_1_548[127:112]   = Conv_out[312];
    assign  image_1_548[111:96]    = Conv_out[311];
    assign  image_1_548[95:80]     = Conv_out[283];
    assign  image_1_548[79:64]     = Conv_out[282];
    assign  image_1_548[63:48]     = Conv_out[281];
    assign  image_1_548[47:32]     = Conv_out[253];
    assign  image_1_548[31:16]     = Conv_out[252];
    assign  image_1_548[15:0]      = Conv_out[251];

    assign  image_1_549[143:128]   = Conv_out[312];
    assign  image_1_549[127:112]   = Conv_out[311];
    assign  image_1_549[111:96]    = Conv_out[310];
    assign  image_1_549[95:80]     = Conv_out[282];
    assign  image_1_549[79:64]     = Conv_out[281];
    assign  image_1_549[63:48]     = Conv_out[280];
    assign  image_1_549[47:32]     = Conv_out[252];
    assign  image_1_549[31:16]     = Conv_out[251];
    assign  image_1_549[15:0]      = Conv_out[250];

    assign  image_1_550[143:128]   = Conv_out[311];
    assign  image_1_550[127:112]   = Conv_out[310];
    assign  image_1_550[111:96]    = Conv_out[309];
    assign  image_1_550[95:80]     = Conv_out[281];
    assign  image_1_550[79:64]     = Conv_out[280];
    assign  image_1_550[63:48]     = Conv_out[279];
    assign  image_1_550[47:32]     = Conv_out[251];
    assign  image_1_550[31:16]     = Conv_out[250];
    assign  image_1_550[15:0]      = Conv_out[249];

    assign  image_1_551[143:128]   = Conv_out[310];
    assign  image_1_551[127:112]   = Conv_out[309];
    assign  image_1_551[111:96]    = Conv_out[308];
    assign  image_1_551[95:80]     = Conv_out[280];
    assign  image_1_551[79:64]     = Conv_out[279];
    assign  image_1_551[63:48]     = Conv_out[278];
    assign  image_1_551[47:32]     = Conv_out[250];
    assign  image_1_551[31:16]     = Conv_out[249];
    assign  image_1_551[15:0]      = Conv_out[248];

    assign  image_1_552[143:128]   = Conv_out[309];
    assign  image_1_552[127:112]   = Conv_out[308];
    assign  image_1_552[111:96]    = Conv_out[307];
    assign  image_1_552[95:80]     = Conv_out[279];
    assign  image_1_552[79:64]     = Conv_out[278];
    assign  image_1_552[63:48]     = Conv_out[277];
    assign  image_1_552[47:32]     = Conv_out[249];
    assign  image_1_552[31:16]     = Conv_out[248];
    assign  image_1_552[15:0]      = Conv_out[247];

    assign  image_1_553[143:128]   = Conv_out[308];
    assign  image_1_553[127:112]   = Conv_out[307];
    assign  image_1_553[111:96]    = Conv_out[306];
    assign  image_1_553[95:80]     = Conv_out[278];
    assign  image_1_553[79:64]     = Conv_out[277];
    assign  image_1_553[63:48]     = Conv_out[276];
    assign  image_1_553[47:32]     = Conv_out[248];
    assign  image_1_553[31:16]     = Conv_out[247];
    assign  image_1_553[15:0]      = Conv_out[246];

    assign  image_1_554[143:128]   = Conv_out[307];
    assign  image_1_554[127:112]   = Conv_out[306];
    assign  image_1_554[111:96]    = Conv_out[305];
    assign  image_1_554[95:80]     = Conv_out[277];
    assign  image_1_554[79:64]     = Conv_out[276];
    assign  image_1_554[63:48]     = Conv_out[275];
    assign  image_1_554[47:32]     = Conv_out[247];
    assign  image_1_554[31:16]     = Conv_out[246];
    assign  image_1_554[15:0]      = Conv_out[245];

    assign  image_1_555[143:128]   = Conv_out[306];
    assign  image_1_555[127:112]   = Conv_out[305];
    assign  image_1_555[111:96]    = Conv_out[304];
    assign  image_1_555[95:80]     = Conv_out[276];
    assign  image_1_555[79:64]     = Conv_out[275];
    assign  image_1_555[63:48]     = Conv_out[274];
    assign  image_1_555[47:32]     = Conv_out[246];
    assign  image_1_555[31:16]     = Conv_out[245];
    assign  image_1_555[15:0]      = Conv_out[244];

    assign  image_1_556[143:128]   = Conv_out[305];
    assign  image_1_556[127:112]   = Conv_out[304];
    assign  image_1_556[111:96]    = Conv_out[303];
    assign  image_1_556[95:80]     = Conv_out[275];
    assign  image_1_556[79:64]     = Conv_out[274];
    assign  image_1_556[63:48]     = Conv_out[273];
    assign  image_1_556[47:32]     = Conv_out[245];
    assign  image_1_556[31:16]     = Conv_out[244];
    assign  image_1_556[15:0]      = Conv_out[243];

    assign  image_1_557[143:128]   = Conv_out[304];
    assign  image_1_557[127:112]   = Conv_out[303];
    assign  image_1_557[111:96]    = Conv_out[302];
    assign  image_1_557[95:80]     = Conv_out[274];
    assign  image_1_557[79:64]     = Conv_out[273];
    assign  image_1_557[63:48]     = Conv_out[272];
    assign  image_1_557[47:32]     = Conv_out[244];
    assign  image_1_557[31:16]     = Conv_out[243];
    assign  image_1_557[15:0]      = Conv_out[242];

    assign  image_1_558[143:128]   = Conv_out[303];
    assign  image_1_558[127:112]   = Conv_out[302];
    assign  image_1_558[111:96]    = Conv_out[301];
    assign  image_1_558[95:80]     = Conv_out[273];
    assign  image_1_558[79:64]     = Conv_out[272];
    assign  image_1_558[63:48]     = Conv_out[271];
    assign  image_1_558[47:32]     = Conv_out[243];
    assign  image_1_558[31:16]     = Conv_out[242];
    assign  image_1_558[15:0]      = Conv_out[241];

    assign  image_1_559[143:128]   = Conv_out[302];
    assign  image_1_559[127:112]   = Conv_out[301];
    assign  image_1_559[111:96]    = Conv_out[300];
    assign  image_1_559[95:80]     = Conv_out[272];
    assign  image_1_559[79:64]     = Conv_out[271];
    assign  image_1_559[63:48]     = Conv_out[270];
    assign  image_1_559[47:32]     = Conv_out[242];
    assign  image_1_559[31:16]     = Conv_out[241];
    assign  image_1_559[15:0]      = Conv_out[240];

    assign  image_1_560[143:128]   = Conv_out[299];
    assign  image_1_560[127:112]   = Conv_out[298];
    assign  image_1_560[111:96]    = Conv_out[297];
    assign  image_1_560[95:80]     = Conv_out[269];
    assign  image_1_560[79:64]     = Conv_out[268];
    assign  image_1_560[63:48]     = Conv_out[267];
    assign  image_1_560[47:32]     = Conv_out[239];
    assign  image_1_560[31:16]     = Conv_out[238];
    assign  image_1_560[15:0]      = Conv_out[237];

    assign  image_1_561[143:128]   = Conv_out[298];
    assign  image_1_561[127:112]   = Conv_out[297];
    assign  image_1_561[111:96]    = Conv_out[296];
    assign  image_1_561[95:80]     = Conv_out[268];
    assign  image_1_561[79:64]     = Conv_out[267];
    assign  image_1_561[63:48]     = Conv_out[266];
    assign  image_1_561[47:32]     = Conv_out[238];
    assign  image_1_561[31:16]     = Conv_out[237];
    assign  image_1_561[15:0]      = Conv_out[236];

    assign  image_1_562[143:128]   = Conv_out[297];
    assign  image_1_562[127:112]   = Conv_out[296];
    assign  image_1_562[111:96]    = Conv_out[295];
    assign  image_1_562[95:80]     = Conv_out[267];
    assign  image_1_562[79:64]     = Conv_out[266];
    assign  image_1_562[63:48]     = Conv_out[265];
    assign  image_1_562[47:32]     = Conv_out[237];
    assign  image_1_562[31:16]     = Conv_out[236];
    assign  image_1_562[15:0]      = Conv_out[235];

    assign  image_1_563[143:128]   = Conv_out[296];
    assign  image_1_563[127:112]   = Conv_out[295];
    assign  image_1_563[111:96]    = Conv_out[294];
    assign  image_1_563[95:80]     = Conv_out[266];
    assign  image_1_563[79:64]     = Conv_out[265];
    assign  image_1_563[63:48]     = Conv_out[264];
    assign  image_1_563[47:32]     = Conv_out[236];
    assign  image_1_563[31:16]     = Conv_out[235];
    assign  image_1_563[15:0]      = Conv_out[234];

    assign  image_1_564[143:128]   = Conv_out[295];
    assign  image_1_564[127:112]   = Conv_out[294];
    assign  image_1_564[111:96]    = Conv_out[293];
    assign  image_1_564[95:80]     = Conv_out[265];
    assign  image_1_564[79:64]     = Conv_out[264];
    assign  image_1_564[63:48]     = Conv_out[263];
    assign  image_1_564[47:32]     = Conv_out[235];
    assign  image_1_564[31:16]     = Conv_out[234];
    assign  image_1_564[15:0]      = Conv_out[233];

    assign  image_1_565[143:128]   = Conv_out[294];
    assign  image_1_565[127:112]   = Conv_out[293];
    assign  image_1_565[111:96]    = Conv_out[292];
    assign  image_1_565[95:80]     = Conv_out[264];
    assign  image_1_565[79:64]     = Conv_out[263];
    assign  image_1_565[63:48]     = Conv_out[262];
    assign  image_1_565[47:32]     = Conv_out[234];
    assign  image_1_565[31:16]     = Conv_out[233];
    assign  image_1_565[15:0]      = Conv_out[232];

    assign  image_1_566[143:128]   = Conv_out[293];
    assign  image_1_566[127:112]   = Conv_out[292];
    assign  image_1_566[111:96]    = Conv_out[291];
    assign  image_1_566[95:80]     = Conv_out[263];
    assign  image_1_566[79:64]     = Conv_out[262];
    assign  image_1_566[63:48]     = Conv_out[261];
    assign  image_1_566[47:32]     = Conv_out[233];
    assign  image_1_566[31:16]     = Conv_out[232];
    assign  image_1_566[15:0]      = Conv_out[231];

    assign  image_1_567[143:128]   = Conv_out[292];
    assign  image_1_567[127:112]   = Conv_out[291];
    assign  image_1_567[111:96]    = Conv_out[290];
    assign  image_1_567[95:80]     = Conv_out[262];
    assign  image_1_567[79:64]     = Conv_out[261];
    assign  image_1_567[63:48]     = Conv_out[260];
    assign  image_1_567[47:32]     = Conv_out[232];
    assign  image_1_567[31:16]     = Conv_out[231];
    assign  image_1_567[15:0]      = Conv_out[230];

    assign  image_1_568[143:128]   = Conv_out[291];
    assign  image_1_568[127:112]   = Conv_out[290];
    assign  image_1_568[111:96]    = Conv_out[289];
    assign  image_1_568[95:80]     = Conv_out[261];
    assign  image_1_568[79:64]     = Conv_out[260];
    assign  image_1_568[63:48]     = Conv_out[259];
    assign  image_1_568[47:32]     = Conv_out[231];
    assign  image_1_568[31:16]     = Conv_out[230];
    assign  image_1_568[15:0]      = Conv_out[229];

    assign  image_1_569[143:128]   = Conv_out[290];
    assign  image_1_569[127:112]   = Conv_out[289];
    assign  image_1_569[111:96]    = Conv_out[288];
    assign  image_1_569[95:80]     = Conv_out[260];
    assign  image_1_569[79:64]     = Conv_out[259];
    assign  image_1_569[63:48]     = Conv_out[258];
    assign  image_1_569[47:32]     = Conv_out[230];
    assign  image_1_569[31:16]     = Conv_out[229];
    assign  image_1_569[15:0]      = Conv_out[228];

    assign  image_1_570[143:128]   = Conv_out[289];
    assign  image_1_570[127:112]   = Conv_out[288];
    assign  image_1_570[111:96]    = Conv_out[287];
    assign  image_1_570[95:80]     = Conv_out[259];
    assign  image_1_570[79:64]     = Conv_out[258];
    assign  image_1_570[63:48]     = Conv_out[257];
    assign  image_1_570[47:32]     = Conv_out[229];
    assign  image_1_570[31:16]     = Conv_out[228];
    assign  image_1_570[15:0]      = Conv_out[227];

    assign  image_1_571[143:128]   = Conv_out[288];
    assign  image_1_571[127:112]   = Conv_out[287];
    assign  image_1_571[111:96]    = Conv_out[286];
    assign  image_1_571[95:80]     = Conv_out[258];
    assign  image_1_571[79:64]     = Conv_out[257];
    assign  image_1_571[63:48]     = Conv_out[256];
    assign  image_1_571[47:32]     = Conv_out[228];
    assign  image_1_571[31:16]     = Conv_out[227];
    assign  image_1_571[15:0]      = Conv_out[226];

    assign  image_1_572[143:128]   = Conv_out[287];
    assign  image_1_572[127:112]   = Conv_out[286];
    assign  image_1_572[111:96]    = Conv_out[285];
    assign  image_1_572[95:80]     = Conv_out[257];
    assign  image_1_572[79:64]     = Conv_out[256];
    assign  image_1_572[63:48]     = Conv_out[255];
    assign  image_1_572[47:32]     = Conv_out[227];
    assign  image_1_572[31:16]     = Conv_out[226];
    assign  image_1_572[15:0]      = Conv_out[225];

    assign  image_1_573[143:128]   = Conv_out[286];
    assign  image_1_573[127:112]   = Conv_out[285];
    assign  image_1_573[111:96]    = Conv_out[284];
    assign  image_1_573[95:80]     = Conv_out[256];
    assign  image_1_573[79:64]     = Conv_out[255];
    assign  image_1_573[63:48]     = Conv_out[254];
    assign  image_1_573[47:32]     = Conv_out[226];
    assign  image_1_573[31:16]     = Conv_out[225];
    assign  image_1_573[15:0]      = Conv_out[224];

    assign  image_1_574[143:128]   = Conv_out[285];
    assign  image_1_574[127:112]   = Conv_out[284];
    assign  image_1_574[111:96]    = Conv_out[283];
    assign  image_1_574[95:80]     = Conv_out[255];
    assign  image_1_574[79:64]     = Conv_out[254];
    assign  image_1_574[63:48]     = Conv_out[253];
    assign  image_1_574[47:32]     = Conv_out[225];
    assign  image_1_574[31:16]     = Conv_out[224];
    assign  image_1_574[15:0]      = Conv_out[223];

    assign  image_1_575[143:128]   = Conv_out[284];
    assign  image_1_575[127:112]   = Conv_out[283];
    assign  image_1_575[111:96]    = Conv_out[282];
    assign  image_1_575[95:80]     = Conv_out[254];
    assign  image_1_575[79:64]     = Conv_out[253];
    assign  image_1_575[63:48]     = Conv_out[252];
    assign  image_1_575[47:32]     = Conv_out[224];
    assign  image_1_575[31:16]     = Conv_out[223];
    assign  image_1_575[15:0]      = Conv_out[222];

    assign  image_1_576[143:128]   = Conv_out[283];
    assign  image_1_576[127:112]   = Conv_out[282];
    assign  image_1_576[111:96]    = Conv_out[281];
    assign  image_1_576[95:80]     = Conv_out[253];
    assign  image_1_576[79:64]     = Conv_out[252];
    assign  image_1_576[63:48]     = Conv_out[251];
    assign  image_1_576[47:32]     = Conv_out[223];
    assign  image_1_576[31:16]     = Conv_out[222];
    assign  image_1_576[15:0]      = Conv_out[221];

    assign  image_1_577[143:128]   = Conv_out[282];
    assign  image_1_577[127:112]   = Conv_out[281];
    assign  image_1_577[111:96]    = Conv_out[280];
    assign  image_1_577[95:80]     = Conv_out[252];
    assign  image_1_577[79:64]     = Conv_out[251];
    assign  image_1_577[63:48]     = Conv_out[250];
    assign  image_1_577[47:32]     = Conv_out[222];
    assign  image_1_577[31:16]     = Conv_out[221];
    assign  image_1_577[15:0]      = Conv_out[220];

    assign  image_1_578[143:128]   = Conv_out[281];
    assign  image_1_578[127:112]   = Conv_out[280];
    assign  image_1_578[111:96]    = Conv_out[279];
    assign  image_1_578[95:80]     = Conv_out[251];
    assign  image_1_578[79:64]     = Conv_out[250];
    assign  image_1_578[63:48]     = Conv_out[249];
    assign  image_1_578[47:32]     = Conv_out[221];
    assign  image_1_578[31:16]     = Conv_out[220];
    assign  image_1_578[15:0]      = Conv_out[219];

    assign  image_1_579[143:128]   = Conv_out[280];
    assign  image_1_579[127:112]   = Conv_out[279];
    assign  image_1_579[111:96]    = Conv_out[278];
    assign  image_1_579[95:80]     = Conv_out[250];
    assign  image_1_579[79:64]     = Conv_out[249];
    assign  image_1_579[63:48]     = Conv_out[248];
    assign  image_1_579[47:32]     = Conv_out[220];
    assign  image_1_579[31:16]     = Conv_out[219];
    assign  image_1_579[15:0]      = Conv_out[218];

    assign  image_1_580[143:128]   = Conv_out[279];
    assign  image_1_580[127:112]   = Conv_out[278];
    assign  image_1_580[111:96]    = Conv_out[277];
    assign  image_1_580[95:80]     = Conv_out[249];
    assign  image_1_580[79:64]     = Conv_out[248];
    assign  image_1_580[63:48]     = Conv_out[247];
    assign  image_1_580[47:32]     = Conv_out[219];
    assign  image_1_580[31:16]     = Conv_out[218];
    assign  image_1_580[15:0]      = Conv_out[217];

    assign  image_1_581[143:128]   = Conv_out[278];
    assign  image_1_581[127:112]   = Conv_out[277];
    assign  image_1_581[111:96]    = Conv_out[276];
    assign  image_1_581[95:80]     = Conv_out[248];
    assign  image_1_581[79:64]     = Conv_out[247];
    assign  image_1_581[63:48]     = Conv_out[246];
    assign  image_1_581[47:32]     = Conv_out[218];
    assign  image_1_581[31:16]     = Conv_out[217];
    assign  image_1_581[15:0]      = Conv_out[216];

    assign  image_1_582[143:128]   = Conv_out[277];
    assign  image_1_582[127:112]   = Conv_out[276];
    assign  image_1_582[111:96]    = Conv_out[275];
    assign  image_1_582[95:80]     = Conv_out[247];
    assign  image_1_582[79:64]     = Conv_out[246];
    assign  image_1_582[63:48]     = Conv_out[245];
    assign  image_1_582[47:32]     = Conv_out[217];
    assign  image_1_582[31:16]     = Conv_out[216];
    assign  image_1_582[15:0]      = Conv_out[215];

    assign  image_1_583[143:128]   = Conv_out[276];
    assign  image_1_583[127:112]   = Conv_out[275];
    assign  image_1_583[111:96]    = Conv_out[274];
    assign  image_1_583[95:80]     = Conv_out[246];
    assign  image_1_583[79:64]     = Conv_out[245];
    assign  image_1_583[63:48]     = Conv_out[244];
    assign  image_1_583[47:32]     = Conv_out[216];
    assign  image_1_583[31:16]     = Conv_out[215];
    assign  image_1_583[15:0]      = Conv_out[214];

    assign  image_1_584[143:128]   = Conv_out[275];
    assign  image_1_584[127:112]   = Conv_out[274];
    assign  image_1_584[111:96]    = Conv_out[273];
    assign  image_1_584[95:80]     = Conv_out[245];
    assign  image_1_584[79:64]     = Conv_out[244];
    assign  image_1_584[63:48]     = Conv_out[243];
    assign  image_1_584[47:32]     = Conv_out[215];
    assign  image_1_584[31:16]     = Conv_out[214];
    assign  image_1_584[15:0]      = Conv_out[213];

    assign  image_1_585[143:128]   = Conv_out[274];
    assign  image_1_585[127:112]   = Conv_out[273];
    assign  image_1_585[111:96]    = Conv_out[272];
    assign  image_1_585[95:80]     = Conv_out[244];
    assign  image_1_585[79:64]     = Conv_out[243];
    assign  image_1_585[63:48]     = Conv_out[242];
    assign  image_1_585[47:32]     = Conv_out[214];
    assign  image_1_585[31:16]     = Conv_out[213];
    assign  image_1_585[15:0]      = Conv_out[212];

    assign  image_1_586[143:128]   = Conv_out[273];
    assign  image_1_586[127:112]   = Conv_out[272];
    assign  image_1_586[111:96]    = Conv_out[271];
    assign  image_1_586[95:80]     = Conv_out[243];
    assign  image_1_586[79:64]     = Conv_out[242];
    assign  image_1_586[63:48]     = Conv_out[241];
    assign  image_1_586[47:32]     = Conv_out[213];
    assign  image_1_586[31:16]     = Conv_out[212];
    assign  image_1_586[15:0]      = Conv_out[211];

    assign  image_1_587[143:128]   = Conv_out[272];
    assign  image_1_587[127:112]   = Conv_out[271];
    assign  image_1_587[111:96]    = Conv_out[270];
    assign  image_1_587[95:80]     = Conv_out[242];
    assign  image_1_587[79:64]     = Conv_out[241];
    assign  image_1_587[63:48]     = Conv_out[240];
    assign  image_1_587[47:32]     = Conv_out[212];
    assign  image_1_587[31:16]     = Conv_out[211];
    assign  image_1_587[15:0]      = Conv_out[210];

    assign  image_1_588[143:128]   = Conv_out[269];
    assign  image_1_588[127:112]   = Conv_out[268];
    assign  image_1_588[111:96]    = Conv_out[267];
    assign  image_1_588[95:80]     = Conv_out[239];
    assign  image_1_588[79:64]     = Conv_out[238];
    assign  image_1_588[63:48]     = Conv_out[237];
    assign  image_1_588[47:32]     = Conv_out[209];
    assign  image_1_588[31:16]     = Conv_out[208];
    assign  image_1_588[15:0]      = Conv_out[207];

    assign  image_1_589[143:128]   = Conv_out[268];
    assign  image_1_589[127:112]   = Conv_out[267];
    assign  image_1_589[111:96]    = Conv_out[266];
    assign  image_1_589[95:80]     = Conv_out[238];
    assign  image_1_589[79:64]     = Conv_out[237];
    assign  image_1_589[63:48]     = Conv_out[236];
    assign  image_1_589[47:32]     = Conv_out[208];
    assign  image_1_589[31:16]     = Conv_out[207];
    assign  image_1_589[15:0]      = Conv_out[206];

    assign  image_1_590[143:128]   = Conv_out[267];
    assign  image_1_590[127:112]   = Conv_out[266];
    assign  image_1_590[111:96]    = Conv_out[265];
    assign  image_1_590[95:80]     = Conv_out[237];
    assign  image_1_590[79:64]     = Conv_out[236];
    assign  image_1_590[63:48]     = Conv_out[235];
    assign  image_1_590[47:32]     = Conv_out[207];
    assign  image_1_590[31:16]     = Conv_out[206];
    assign  image_1_590[15:0]      = Conv_out[205];

    assign  image_1_591[143:128]   = Conv_out[266];
    assign  image_1_591[127:112]   = Conv_out[265];
    assign  image_1_591[111:96]    = Conv_out[264];
    assign  image_1_591[95:80]     = Conv_out[236];
    assign  image_1_591[79:64]     = Conv_out[235];
    assign  image_1_591[63:48]     = Conv_out[234];
    assign  image_1_591[47:32]     = Conv_out[206];
    assign  image_1_591[31:16]     = Conv_out[205];
    assign  image_1_591[15:0]      = Conv_out[204];

    assign  image_1_592[143:128]   = Conv_out[265];
    assign  image_1_592[127:112]   = Conv_out[264];
    assign  image_1_592[111:96]    = Conv_out[263];
    assign  image_1_592[95:80]     = Conv_out[235];
    assign  image_1_592[79:64]     = Conv_out[234];
    assign  image_1_592[63:48]     = Conv_out[233];
    assign  image_1_592[47:32]     = Conv_out[205];
    assign  image_1_592[31:16]     = Conv_out[204];
    assign  image_1_592[15:0]      = Conv_out[203];

    assign  image_1_593[143:128]   = Conv_out[264];
    assign  image_1_593[127:112]   = Conv_out[263];
    assign  image_1_593[111:96]    = Conv_out[262];
    assign  image_1_593[95:80]     = Conv_out[234];
    assign  image_1_593[79:64]     = Conv_out[233];
    assign  image_1_593[63:48]     = Conv_out[232];
    assign  image_1_593[47:32]     = Conv_out[204];
    assign  image_1_593[31:16]     = Conv_out[203];
    assign  image_1_593[15:0]      = Conv_out[202];

    assign  image_1_594[143:128]   = Conv_out[263];
    assign  image_1_594[127:112]   = Conv_out[262];
    assign  image_1_594[111:96]    = Conv_out[261];
    assign  image_1_594[95:80]     = Conv_out[233];
    assign  image_1_594[79:64]     = Conv_out[232];
    assign  image_1_594[63:48]     = Conv_out[231];
    assign  image_1_594[47:32]     = Conv_out[203];
    assign  image_1_594[31:16]     = Conv_out[202];
    assign  image_1_594[15:0]      = Conv_out[201];

    assign  image_1_595[143:128]   = Conv_out[262];
    assign  image_1_595[127:112]   = Conv_out[261];
    assign  image_1_595[111:96]    = Conv_out[260];
    assign  image_1_595[95:80]     = Conv_out[232];
    assign  image_1_595[79:64]     = Conv_out[231];
    assign  image_1_595[63:48]     = Conv_out[230];
    assign  image_1_595[47:32]     = Conv_out[202];
    assign  image_1_595[31:16]     = Conv_out[201];
    assign  image_1_595[15:0]      = Conv_out[200];

    assign  image_1_596[143:128]   = Conv_out[261];
    assign  image_1_596[127:112]   = Conv_out[260];
    assign  image_1_596[111:96]    = Conv_out[259];
    assign  image_1_596[95:80]     = Conv_out[231];
    assign  image_1_596[79:64]     = Conv_out[230];
    assign  image_1_596[63:48]     = Conv_out[229];
    assign  image_1_596[47:32]     = Conv_out[201];
    assign  image_1_596[31:16]     = Conv_out[200];
    assign  image_1_596[15:0]      = Conv_out[199];

    assign  image_1_597[143:128]   = Conv_out[260];
    assign  image_1_597[127:112]   = Conv_out[259];
    assign  image_1_597[111:96]    = Conv_out[258];
    assign  image_1_597[95:80]     = Conv_out[230];
    assign  image_1_597[79:64]     = Conv_out[229];
    assign  image_1_597[63:48]     = Conv_out[228];
    assign  image_1_597[47:32]     = Conv_out[200];
    assign  image_1_597[31:16]     = Conv_out[199];
    assign  image_1_597[15:0]      = Conv_out[198];

    assign  image_1_598[143:128]   = Conv_out[259];
    assign  image_1_598[127:112]   = Conv_out[258];
    assign  image_1_598[111:96]    = Conv_out[257];
    assign  image_1_598[95:80]     = Conv_out[229];
    assign  image_1_598[79:64]     = Conv_out[228];
    assign  image_1_598[63:48]     = Conv_out[227];
    assign  image_1_598[47:32]     = Conv_out[199];
    assign  image_1_598[31:16]     = Conv_out[198];
    assign  image_1_598[15:0]      = Conv_out[197];

    assign  image_1_599[143:128]   = Conv_out[258];
    assign  image_1_599[127:112]   = Conv_out[257];
    assign  image_1_599[111:96]    = Conv_out[256];
    assign  image_1_599[95:80]     = Conv_out[228];
    assign  image_1_599[79:64]     = Conv_out[227];
    assign  image_1_599[63:48]     = Conv_out[226];
    assign  image_1_599[47:32]     = Conv_out[198];
    assign  image_1_599[31:16]     = Conv_out[197];
    assign  image_1_599[15:0]      = Conv_out[196];

    assign  image_1_600[143:128]   = Conv_out[257];
    assign  image_1_600[127:112]   = Conv_out[256];
    assign  image_1_600[111:96]    = Conv_out[255];
    assign  image_1_600[95:80]     = Conv_out[227];
    assign  image_1_600[79:64]     = Conv_out[226];
    assign  image_1_600[63:48]     = Conv_out[225];
    assign  image_1_600[47:32]     = Conv_out[197];
    assign  image_1_600[31:16]     = Conv_out[196];
    assign  image_1_600[15:0]      = Conv_out[195];

    assign  image_1_601[143:128]   = Conv_out[256];
    assign  image_1_601[127:112]   = Conv_out[255];
    assign  image_1_601[111:96]    = Conv_out[254];
    assign  image_1_601[95:80]     = Conv_out[226];
    assign  image_1_601[79:64]     = Conv_out[225];
    assign  image_1_601[63:48]     = Conv_out[224];
    assign  image_1_601[47:32]     = Conv_out[196];
    assign  image_1_601[31:16]     = Conv_out[195];
    assign  image_1_601[15:0]      = Conv_out[194];

    assign  image_1_602[143:128]   = Conv_out[255];
    assign  image_1_602[127:112]   = Conv_out[254];
    assign  image_1_602[111:96]    = Conv_out[253];
    assign  image_1_602[95:80]     = Conv_out[225];
    assign  image_1_602[79:64]     = Conv_out[224];
    assign  image_1_602[63:48]     = Conv_out[223];
    assign  image_1_602[47:32]     = Conv_out[195];
    assign  image_1_602[31:16]     = Conv_out[194];
    assign  image_1_602[15:0]      = Conv_out[193];

    assign  image_1_603[143:128]   = Conv_out[254];
    assign  image_1_603[127:112]   = Conv_out[253];
    assign  image_1_603[111:96]    = Conv_out[252];
    assign  image_1_603[95:80]     = Conv_out[224];
    assign  image_1_603[79:64]     = Conv_out[223];
    assign  image_1_603[63:48]     = Conv_out[222];
    assign  image_1_603[47:32]     = Conv_out[194];
    assign  image_1_603[31:16]     = Conv_out[193];
    assign  image_1_603[15:0]      = Conv_out[192];

    assign  image_1_604[143:128]   = Conv_out[253];
    assign  image_1_604[127:112]   = Conv_out[252];
    assign  image_1_604[111:96]    = Conv_out[251];
    assign  image_1_604[95:80]     = Conv_out[223];
    assign  image_1_604[79:64]     = Conv_out[222];
    assign  image_1_604[63:48]     = Conv_out[221];
    assign  image_1_604[47:32]     = Conv_out[193];
    assign  image_1_604[31:16]     = Conv_out[192];
    assign  image_1_604[15:0]      = Conv_out[191];

    assign  image_1_605[143:128]   = Conv_out[252];
    assign  image_1_605[127:112]   = Conv_out[251];
    assign  image_1_605[111:96]    = Conv_out[250];
    assign  image_1_605[95:80]     = Conv_out[222];
    assign  image_1_605[79:64]     = Conv_out[221];
    assign  image_1_605[63:48]     = Conv_out[220];
    assign  image_1_605[47:32]     = Conv_out[192];
    assign  image_1_605[31:16]     = Conv_out[191];
    assign  image_1_605[15:0]      = Conv_out[190];

    assign  image_1_606[143:128]   = Conv_out[251];
    assign  image_1_606[127:112]   = Conv_out[250];
    assign  image_1_606[111:96]    = Conv_out[249];
    assign  image_1_606[95:80]     = Conv_out[221];
    assign  image_1_606[79:64]     = Conv_out[220];
    assign  image_1_606[63:48]     = Conv_out[219];
    assign  image_1_606[47:32]     = Conv_out[191];
    assign  image_1_606[31:16]     = Conv_out[190];
    assign  image_1_606[15:0]      = Conv_out[189];

    assign  image_1_607[143:128]   = Conv_out[250];
    assign  image_1_607[127:112]   = Conv_out[249];
    assign  image_1_607[111:96]    = Conv_out[248];
    assign  image_1_607[95:80]     = Conv_out[220];
    assign  image_1_607[79:64]     = Conv_out[219];
    assign  image_1_607[63:48]     = Conv_out[218];
    assign  image_1_607[47:32]     = Conv_out[190];
    assign  image_1_607[31:16]     = Conv_out[189];
    assign  image_1_607[15:0]      = Conv_out[188];

    assign  image_1_608[143:128]   = Conv_out[249];
    assign  image_1_608[127:112]   = Conv_out[248];
    assign  image_1_608[111:96]    = Conv_out[247];
    assign  image_1_608[95:80]     = Conv_out[219];
    assign  image_1_608[79:64]     = Conv_out[218];
    assign  image_1_608[63:48]     = Conv_out[217];
    assign  image_1_608[47:32]     = Conv_out[189];
    assign  image_1_608[31:16]     = Conv_out[188];
    assign  image_1_608[15:0]      = Conv_out[187];

    assign  image_1_609[143:128]   = Conv_out[248];
    assign  image_1_609[127:112]   = Conv_out[247];
    assign  image_1_609[111:96]    = Conv_out[246];
    assign  image_1_609[95:80]     = Conv_out[218];
    assign  image_1_609[79:64]     = Conv_out[217];
    assign  image_1_609[63:48]     = Conv_out[216];
    assign  image_1_609[47:32]     = Conv_out[188];
    assign  image_1_609[31:16]     = Conv_out[187];
    assign  image_1_609[15:0]      = Conv_out[186];

    assign  image_1_610[143:128]   = Conv_out[247];
    assign  image_1_610[127:112]   = Conv_out[246];
    assign  image_1_610[111:96]    = Conv_out[245];
    assign  image_1_610[95:80]     = Conv_out[217];
    assign  image_1_610[79:64]     = Conv_out[216];
    assign  image_1_610[63:48]     = Conv_out[215];
    assign  image_1_610[47:32]     = Conv_out[187];
    assign  image_1_610[31:16]     = Conv_out[186];
    assign  image_1_610[15:0]      = Conv_out[185];

    assign  image_1_611[143:128]   = Conv_out[246];
    assign  image_1_611[127:112]   = Conv_out[245];
    assign  image_1_611[111:96]    = Conv_out[244];
    assign  image_1_611[95:80]     = Conv_out[216];
    assign  image_1_611[79:64]     = Conv_out[215];
    assign  image_1_611[63:48]     = Conv_out[214];
    assign  image_1_611[47:32]     = Conv_out[186];
    assign  image_1_611[31:16]     = Conv_out[185];
    assign  image_1_611[15:0]      = Conv_out[184];

    assign  image_1_612[143:128]   = Conv_out[245];
    assign  image_1_612[127:112]   = Conv_out[244];
    assign  image_1_612[111:96]    = Conv_out[243];
    assign  image_1_612[95:80]     = Conv_out[215];
    assign  image_1_612[79:64]     = Conv_out[214];
    assign  image_1_612[63:48]     = Conv_out[213];
    assign  image_1_612[47:32]     = Conv_out[185];
    assign  image_1_612[31:16]     = Conv_out[184];
    assign  image_1_612[15:0]      = Conv_out[183];

    assign  image_1_613[143:128]   = Conv_out[244];
    assign  image_1_613[127:112]   = Conv_out[243];
    assign  image_1_613[111:96]    = Conv_out[242];
    assign  image_1_613[95:80]     = Conv_out[214];
    assign  image_1_613[79:64]     = Conv_out[213];
    assign  image_1_613[63:48]     = Conv_out[212];
    assign  image_1_613[47:32]     = Conv_out[184];
    assign  image_1_613[31:16]     = Conv_out[183];
    assign  image_1_613[15:0]      = Conv_out[182];

    assign  image_1_614[143:128]   = Conv_out[243];
    assign  image_1_614[127:112]   = Conv_out[242];
    assign  image_1_614[111:96]    = Conv_out[241];
    assign  image_1_614[95:80]     = Conv_out[213];
    assign  image_1_614[79:64]     = Conv_out[212];
    assign  image_1_614[63:48]     = Conv_out[211];
    assign  image_1_614[47:32]     = Conv_out[183];
    assign  image_1_614[31:16]     = Conv_out[182];
    assign  image_1_614[15:0]      = Conv_out[181];

    assign  image_1_615[143:128]   = Conv_out[242];
    assign  image_1_615[127:112]   = Conv_out[241];
    assign  image_1_615[111:96]    = Conv_out[240];
    assign  image_1_615[95:80]     = Conv_out[212];
    assign  image_1_615[79:64]     = Conv_out[211];
    assign  image_1_615[63:48]     = Conv_out[210];
    assign  image_1_615[47:32]     = Conv_out[182];
    assign  image_1_615[31:16]     = Conv_out[181];
    assign  image_1_615[15:0]      = Conv_out[180];

    assign  image_1_616[143:128]   = Conv_out[239];
    assign  image_1_616[127:112]   = Conv_out[238];
    assign  image_1_616[111:96]    = Conv_out[237];
    assign  image_1_616[95:80]     = Conv_out[209];
    assign  image_1_616[79:64]     = Conv_out[208];
    assign  image_1_616[63:48]     = Conv_out[207];
    assign  image_1_616[47:32]     = Conv_out[179];
    assign  image_1_616[31:16]     = Conv_out[178];
    assign  image_1_616[15:0]      = Conv_out[177];

    assign  image_1_617[143:128]   = Conv_out[238];
    assign  image_1_617[127:112]   = Conv_out[237];
    assign  image_1_617[111:96]    = Conv_out[236];
    assign  image_1_617[95:80]     = Conv_out[208];
    assign  image_1_617[79:64]     = Conv_out[207];
    assign  image_1_617[63:48]     = Conv_out[206];
    assign  image_1_617[47:32]     = Conv_out[178];
    assign  image_1_617[31:16]     = Conv_out[177];
    assign  image_1_617[15:0]      = Conv_out[176];

    assign  image_1_618[143:128]   = Conv_out[237];
    assign  image_1_618[127:112]   = Conv_out[236];
    assign  image_1_618[111:96]    = Conv_out[235];
    assign  image_1_618[95:80]     = Conv_out[207];
    assign  image_1_618[79:64]     = Conv_out[206];
    assign  image_1_618[63:48]     = Conv_out[205];
    assign  image_1_618[47:32]     = Conv_out[177];
    assign  image_1_618[31:16]     = Conv_out[176];
    assign  image_1_618[15:0]      = Conv_out[175];

    assign  image_1_619[143:128]   = Conv_out[236];
    assign  image_1_619[127:112]   = Conv_out[235];
    assign  image_1_619[111:96]    = Conv_out[234];
    assign  image_1_619[95:80]     = Conv_out[206];
    assign  image_1_619[79:64]     = Conv_out[205];
    assign  image_1_619[63:48]     = Conv_out[204];
    assign  image_1_619[47:32]     = Conv_out[176];
    assign  image_1_619[31:16]     = Conv_out[175];
    assign  image_1_619[15:0]      = Conv_out[174];

    assign  image_1_620[143:128]   = Conv_out[235];
    assign  image_1_620[127:112]   = Conv_out[234];
    assign  image_1_620[111:96]    = Conv_out[233];
    assign  image_1_620[95:80]     = Conv_out[205];
    assign  image_1_620[79:64]     = Conv_out[204];
    assign  image_1_620[63:48]     = Conv_out[203];
    assign  image_1_620[47:32]     = Conv_out[175];
    assign  image_1_620[31:16]     = Conv_out[174];
    assign  image_1_620[15:0]      = Conv_out[173];

    assign  image_1_621[143:128]   = Conv_out[234];
    assign  image_1_621[127:112]   = Conv_out[233];
    assign  image_1_621[111:96]    = Conv_out[232];
    assign  image_1_621[95:80]     = Conv_out[204];
    assign  image_1_621[79:64]     = Conv_out[203];
    assign  image_1_621[63:48]     = Conv_out[202];
    assign  image_1_621[47:32]     = Conv_out[174];
    assign  image_1_621[31:16]     = Conv_out[173];
    assign  image_1_621[15:0]      = Conv_out[172];

    assign  image_1_622[143:128]   = Conv_out[233];
    assign  image_1_622[127:112]   = Conv_out[232];
    assign  image_1_622[111:96]    = Conv_out[231];
    assign  image_1_622[95:80]     = Conv_out[203];
    assign  image_1_622[79:64]     = Conv_out[202];
    assign  image_1_622[63:48]     = Conv_out[201];
    assign  image_1_622[47:32]     = Conv_out[173];
    assign  image_1_622[31:16]     = Conv_out[172];
    assign  image_1_622[15:0]      = Conv_out[171];

    assign  image_1_623[143:128]   = Conv_out[232];
    assign  image_1_623[127:112]   = Conv_out[231];
    assign  image_1_623[111:96]    = Conv_out[230];
    assign  image_1_623[95:80]     = Conv_out[202];
    assign  image_1_623[79:64]     = Conv_out[201];
    assign  image_1_623[63:48]     = Conv_out[200];
    assign  image_1_623[47:32]     = Conv_out[172];
    assign  image_1_623[31:16]     = Conv_out[171];
    assign  image_1_623[15:0]      = Conv_out[170];

    assign  image_1_624[143:128]   = Conv_out[231];
    assign  image_1_624[127:112]   = Conv_out[230];
    assign  image_1_624[111:96]    = Conv_out[229];
    assign  image_1_624[95:80]     = Conv_out[201];
    assign  image_1_624[79:64]     = Conv_out[200];
    assign  image_1_624[63:48]     = Conv_out[199];
    assign  image_1_624[47:32]     = Conv_out[171];
    assign  image_1_624[31:16]     = Conv_out[170];
    assign  image_1_624[15:0]      = Conv_out[169];

    assign  image_1_625[143:128]   = Conv_out[230];
    assign  image_1_625[127:112]   = Conv_out[229];
    assign  image_1_625[111:96]    = Conv_out[228];
    assign  image_1_625[95:80]     = Conv_out[200];
    assign  image_1_625[79:64]     = Conv_out[199];
    assign  image_1_625[63:48]     = Conv_out[198];
    assign  image_1_625[47:32]     = Conv_out[170];
    assign  image_1_625[31:16]     = Conv_out[169];
    assign  image_1_625[15:0]      = Conv_out[168];

    assign  image_1_626[143:128]   = Conv_out[229];
    assign  image_1_626[127:112]   = Conv_out[228];
    assign  image_1_626[111:96]    = Conv_out[227];
    assign  image_1_626[95:80]     = Conv_out[199];
    assign  image_1_626[79:64]     = Conv_out[198];
    assign  image_1_626[63:48]     = Conv_out[197];
    assign  image_1_626[47:32]     = Conv_out[169];
    assign  image_1_626[31:16]     = Conv_out[168];
    assign  image_1_626[15:0]      = Conv_out[167];

    assign  image_1_627[143:128]   = Conv_out[228];
    assign  image_1_627[127:112]   = Conv_out[227];
    assign  image_1_627[111:96]    = Conv_out[226];
    assign  image_1_627[95:80]     = Conv_out[198];
    assign  image_1_627[79:64]     = Conv_out[197];
    assign  image_1_627[63:48]     = Conv_out[196];
    assign  image_1_627[47:32]     = Conv_out[168];
    assign  image_1_627[31:16]     = Conv_out[167];
    assign  image_1_627[15:0]      = Conv_out[166];

    assign  image_1_628[143:128]   = Conv_out[227];
    assign  image_1_628[127:112]   = Conv_out[226];
    assign  image_1_628[111:96]    = Conv_out[225];
    assign  image_1_628[95:80]     = Conv_out[197];
    assign  image_1_628[79:64]     = Conv_out[196];
    assign  image_1_628[63:48]     = Conv_out[195];
    assign  image_1_628[47:32]     = Conv_out[167];
    assign  image_1_628[31:16]     = Conv_out[166];
    assign  image_1_628[15:0]      = Conv_out[165];

    assign  image_1_629[143:128]   = Conv_out[226];
    assign  image_1_629[127:112]   = Conv_out[225];
    assign  image_1_629[111:96]    = Conv_out[224];
    assign  image_1_629[95:80]     = Conv_out[196];
    assign  image_1_629[79:64]     = Conv_out[195];
    assign  image_1_629[63:48]     = Conv_out[194];
    assign  image_1_629[47:32]     = Conv_out[166];
    assign  image_1_629[31:16]     = Conv_out[165];
    assign  image_1_629[15:0]      = Conv_out[164];

    assign  image_1_630[143:128]   = Conv_out[225];
    assign  image_1_630[127:112]   = Conv_out[224];
    assign  image_1_630[111:96]    = Conv_out[223];
    assign  image_1_630[95:80]     = Conv_out[195];
    assign  image_1_630[79:64]     = Conv_out[194];
    assign  image_1_630[63:48]     = Conv_out[193];
    assign  image_1_630[47:32]     = Conv_out[165];
    assign  image_1_630[31:16]     = Conv_out[164];
    assign  image_1_630[15:0]      = Conv_out[163];

    assign  image_1_631[143:128]   = Conv_out[224];
    assign  image_1_631[127:112]   = Conv_out[223];
    assign  image_1_631[111:96]    = Conv_out[222];
    assign  image_1_631[95:80]     = Conv_out[194];
    assign  image_1_631[79:64]     = Conv_out[193];
    assign  image_1_631[63:48]     = Conv_out[192];
    assign  image_1_631[47:32]     = Conv_out[164];
    assign  image_1_631[31:16]     = Conv_out[163];
    assign  image_1_631[15:0]      = Conv_out[162];

    assign  image_1_632[143:128]   = Conv_out[223];
    assign  image_1_632[127:112]   = Conv_out[222];
    assign  image_1_632[111:96]    = Conv_out[221];
    assign  image_1_632[95:80]     = Conv_out[193];
    assign  image_1_632[79:64]     = Conv_out[192];
    assign  image_1_632[63:48]     = Conv_out[191];
    assign  image_1_632[47:32]     = Conv_out[163];
    assign  image_1_632[31:16]     = Conv_out[162];
    assign  image_1_632[15:0]      = Conv_out[161];

    assign  image_1_633[143:128]   = Conv_out[222];
    assign  image_1_633[127:112]   = Conv_out[221];
    assign  image_1_633[111:96]    = Conv_out[220];
    assign  image_1_633[95:80]     = Conv_out[192];
    assign  image_1_633[79:64]     = Conv_out[191];
    assign  image_1_633[63:48]     = Conv_out[190];
    assign  image_1_633[47:32]     = Conv_out[162];
    assign  image_1_633[31:16]     = Conv_out[161];
    assign  image_1_633[15:0]      = Conv_out[160];

    assign  image_1_634[143:128]   = Conv_out[221];
    assign  image_1_634[127:112]   = Conv_out[220];
    assign  image_1_634[111:96]    = Conv_out[219];
    assign  image_1_634[95:80]     = Conv_out[191];
    assign  image_1_634[79:64]     = Conv_out[190];
    assign  image_1_634[63:48]     = Conv_out[189];
    assign  image_1_634[47:32]     = Conv_out[161];
    assign  image_1_634[31:16]     = Conv_out[160];
    assign  image_1_634[15:0]      = Conv_out[159];

    assign  image_1_635[143:128]   = Conv_out[220];
    assign  image_1_635[127:112]   = Conv_out[219];
    assign  image_1_635[111:96]    = Conv_out[218];
    assign  image_1_635[95:80]     = Conv_out[190];
    assign  image_1_635[79:64]     = Conv_out[189];
    assign  image_1_635[63:48]     = Conv_out[188];
    assign  image_1_635[47:32]     = Conv_out[160];
    assign  image_1_635[31:16]     = Conv_out[159];
    assign  image_1_635[15:0]      = Conv_out[158];

    assign  image_1_636[143:128]   = Conv_out[219];
    assign  image_1_636[127:112]   = Conv_out[218];
    assign  image_1_636[111:96]    = Conv_out[217];
    assign  image_1_636[95:80]     = Conv_out[189];
    assign  image_1_636[79:64]     = Conv_out[188];
    assign  image_1_636[63:48]     = Conv_out[187];
    assign  image_1_636[47:32]     = Conv_out[159];
    assign  image_1_636[31:16]     = Conv_out[158];
    assign  image_1_636[15:0]      = Conv_out[157];

    assign  image_1_637[143:128]   = Conv_out[218];
    assign  image_1_637[127:112]   = Conv_out[217];
    assign  image_1_637[111:96]    = Conv_out[216];
    assign  image_1_637[95:80]     = Conv_out[188];
    assign  image_1_637[79:64]     = Conv_out[187];
    assign  image_1_637[63:48]     = Conv_out[186];
    assign  image_1_637[47:32]     = Conv_out[158];
    assign  image_1_637[31:16]     = Conv_out[157];
    assign  image_1_637[15:0]      = Conv_out[156];

    assign  image_1_638[143:128]   = Conv_out[217];
    assign  image_1_638[127:112]   = Conv_out[216];
    assign  image_1_638[111:96]    = Conv_out[215];
    assign  image_1_638[95:80]     = Conv_out[187];
    assign  image_1_638[79:64]     = Conv_out[186];
    assign  image_1_638[63:48]     = Conv_out[185];
    assign  image_1_638[47:32]     = Conv_out[157];
    assign  image_1_638[31:16]     = Conv_out[156];
    assign  image_1_638[15:0]      = Conv_out[155];

    assign  image_1_639[143:128]   = Conv_out[216];
    assign  image_1_639[127:112]   = Conv_out[215];
    assign  image_1_639[111:96]    = Conv_out[214];
    assign  image_1_639[95:80]     = Conv_out[186];
    assign  image_1_639[79:64]     = Conv_out[185];
    assign  image_1_639[63:48]     = Conv_out[184];
    assign  image_1_639[47:32]     = Conv_out[156];
    assign  image_1_639[31:16]     = Conv_out[155];
    assign  image_1_639[15:0]      = Conv_out[154];

    assign  image_1_640[143:128]   = Conv_out[215];
    assign  image_1_640[127:112]   = Conv_out[214];
    assign  image_1_640[111:96]    = Conv_out[213];
    assign  image_1_640[95:80]     = Conv_out[185];
    assign  image_1_640[79:64]     = Conv_out[184];
    assign  image_1_640[63:48]     = Conv_out[183];
    assign  image_1_640[47:32]     = Conv_out[155];
    assign  image_1_640[31:16]     = Conv_out[154];
    assign  image_1_640[15:0]      = Conv_out[153];

    assign  image_1_641[143:128]   = Conv_out[214];
    assign  image_1_641[127:112]   = Conv_out[213];
    assign  image_1_641[111:96]    = Conv_out[212];
    assign  image_1_641[95:80]     = Conv_out[184];
    assign  image_1_641[79:64]     = Conv_out[183];
    assign  image_1_641[63:48]     = Conv_out[182];
    assign  image_1_641[47:32]     = Conv_out[154];
    assign  image_1_641[31:16]     = Conv_out[153];
    assign  image_1_641[15:0]      = Conv_out[152];

    assign  image_1_642[143:128]   = Conv_out[213];
    assign  image_1_642[127:112]   = Conv_out[212];
    assign  image_1_642[111:96]    = Conv_out[211];
    assign  image_1_642[95:80]     = Conv_out[183];
    assign  image_1_642[79:64]     = Conv_out[182];
    assign  image_1_642[63:48]     = Conv_out[181];
    assign  image_1_642[47:32]     = Conv_out[153];
    assign  image_1_642[31:16]     = Conv_out[152];
    assign  image_1_642[15:0]      = Conv_out[151];

    assign  image_1_643[143:128]   = Conv_out[212];
    assign  image_1_643[127:112]   = Conv_out[211];
    assign  image_1_643[111:96]    = Conv_out[210];
    assign  image_1_643[95:80]     = Conv_out[182];
    assign  image_1_643[79:64]     = Conv_out[181];
    assign  image_1_643[63:48]     = Conv_out[180];
    assign  image_1_643[47:32]     = Conv_out[152];
    assign  image_1_643[31:16]     = Conv_out[151];
    assign  image_1_643[15:0]      = Conv_out[150];

    assign  image_1_644[143:128]   = Conv_out[209];
    assign  image_1_644[127:112]   = Conv_out[208];
    assign  image_1_644[111:96]    = Conv_out[207];
    assign  image_1_644[95:80]     = Conv_out[179];
    assign  image_1_644[79:64]     = Conv_out[178];
    assign  image_1_644[63:48]     = Conv_out[177];
    assign  image_1_644[47:32]     = Conv_out[149];
    assign  image_1_644[31:16]     = Conv_out[148];
    assign  image_1_644[15:0]      = Conv_out[147];

    assign  image_1_645[143:128]   = Conv_out[208];
    assign  image_1_645[127:112]   = Conv_out[207];
    assign  image_1_645[111:96]    = Conv_out[206];
    assign  image_1_645[95:80]     = Conv_out[178];
    assign  image_1_645[79:64]     = Conv_out[177];
    assign  image_1_645[63:48]     = Conv_out[176];
    assign  image_1_645[47:32]     = Conv_out[148];
    assign  image_1_645[31:16]     = Conv_out[147];
    assign  image_1_645[15:0]      = Conv_out[146];

    assign  image_1_646[143:128]   = Conv_out[207];
    assign  image_1_646[127:112]   = Conv_out[206];
    assign  image_1_646[111:96]    = Conv_out[205];
    assign  image_1_646[95:80]     = Conv_out[177];
    assign  image_1_646[79:64]     = Conv_out[176];
    assign  image_1_646[63:48]     = Conv_out[175];
    assign  image_1_646[47:32]     = Conv_out[147];
    assign  image_1_646[31:16]     = Conv_out[146];
    assign  image_1_646[15:0]      = Conv_out[145];

    assign  image_1_647[143:128]   = Conv_out[206];
    assign  image_1_647[127:112]   = Conv_out[205];
    assign  image_1_647[111:96]    = Conv_out[204];
    assign  image_1_647[95:80]     = Conv_out[176];
    assign  image_1_647[79:64]     = Conv_out[175];
    assign  image_1_647[63:48]     = Conv_out[174];
    assign  image_1_647[47:32]     = Conv_out[146];
    assign  image_1_647[31:16]     = Conv_out[145];
    assign  image_1_647[15:0]      = Conv_out[144];

    assign  image_1_648[143:128]   = Conv_out[205];
    assign  image_1_648[127:112]   = Conv_out[204];
    assign  image_1_648[111:96]    = Conv_out[203];
    assign  image_1_648[95:80]     = Conv_out[175];
    assign  image_1_648[79:64]     = Conv_out[174];
    assign  image_1_648[63:48]     = Conv_out[173];
    assign  image_1_648[47:32]     = Conv_out[145];
    assign  image_1_648[31:16]     = Conv_out[144];
    assign  image_1_648[15:0]      = Conv_out[143];

    assign  image_1_649[143:128]   = Conv_out[204];
    assign  image_1_649[127:112]   = Conv_out[203];
    assign  image_1_649[111:96]    = Conv_out[202];
    assign  image_1_649[95:80]     = Conv_out[174];
    assign  image_1_649[79:64]     = Conv_out[173];
    assign  image_1_649[63:48]     = Conv_out[172];
    assign  image_1_649[47:32]     = Conv_out[144];
    assign  image_1_649[31:16]     = Conv_out[143];
    assign  image_1_649[15:0]      = Conv_out[142];

    assign  image_1_650[143:128]   = Conv_out[203];
    assign  image_1_650[127:112]   = Conv_out[202];
    assign  image_1_650[111:96]    = Conv_out[201];
    assign  image_1_650[95:80]     = Conv_out[173];
    assign  image_1_650[79:64]     = Conv_out[172];
    assign  image_1_650[63:48]     = Conv_out[171];
    assign  image_1_650[47:32]     = Conv_out[143];
    assign  image_1_650[31:16]     = Conv_out[142];
    assign  image_1_650[15:0]      = Conv_out[141];

    assign  image_1_651[143:128]   = Conv_out[202];
    assign  image_1_651[127:112]   = Conv_out[201];
    assign  image_1_651[111:96]    = Conv_out[200];
    assign  image_1_651[95:80]     = Conv_out[172];
    assign  image_1_651[79:64]     = Conv_out[171];
    assign  image_1_651[63:48]     = Conv_out[170];
    assign  image_1_651[47:32]     = Conv_out[142];
    assign  image_1_651[31:16]     = Conv_out[141];
    assign  image_1_651[15:0]      = Conv_out[140];

    assign  image_1_652[143:128]   = Conv_out[201];
    assign  image_1_652[127:112]   = Conv_out[200];
    assign  image_1_652[111:96]    = Conv_out[199];
    assign  image_1_652[95:80]     = Conv_out[171];
    assign  image_1_652[79:64]     = Conv_out[170];
    assign  image_1_652[63:48]     = Conv_out[169];
    assign  image_1_652[47:32]     = Conv_out[141];
    assign  image_1_652[31:16]     = Conv_out[140];
    assign  image_1_652[15:0]      = Conv_out[139];

    assign  image_1_653[143:128]   = Conv_out[200];
    assign  image_1_653[127:112]   = Conv_out[199];
    assign  image_1_653[111:96]    = Conv_out[198];
    assign  image_1_653[95:80]     = Conv_out[170];
    assign  image_1_653[79:64]     = Conv_out[169];
    assign  image_1_653[63:48]     = Conv_out[168];
    assign  image_1_653[47:32]     = Conv_out[140];
    assign  image_1_653[31:16]     = Conv_out[139];
    assign  image_1_653[15:0]      = Conv_out[138];

    assign  image_1_654[143:128]   = Conv_out[199];
    assign  image_1_654[127:112]   = Conv_out[198];
    assign  image_1_654[111:96]    = Conv_out[197];
    assign  image_1_654[95:80]     = Conv_out[169];
    assign  image_1_654[79:64]     = Conv_out[168];
    assign  image_1_654[63:48]     = Conv_out[167];
    assign  image_1_654[47:32]     = Conv_out[139];
    assign  image_1_654[31:16]     = Conv_out[138];
    assign  image_1_654[15:0]      = Conv_out[137];

    assign  image_1_655[143:128]   = Conv_out[198];
    assign  image_1_655[127:112]   = Conv_out[197];
    assign  image_1_655[111:96]    = Conv_out[196];
    assign  image_1_655[95:80]     = Conv_out[168];
    assign  image_1_655[79:64]     = Conv_out[167];
    assign  image_1_655[63:48]     = Conv_out[166];
    assign  image_1_655[47:32]     = Conv_out[138];
    assign  image_1_655[31:16]     = Conv_out[137];
    assign  image_1_655[15:0]      = Conv_out[136];

    assign  image_1_656[143:128]   = Conv_out[197];
    assign  image_1_656[127:112]   = Conv_out[196];
    assign  image_1_656[111:96]    = Conv_out[195];
    assign  image_1_656[95:80]     = Conv_out[167];
    assign  image_1_656[79:64]     = Conv_out[166];
    assign  image_1_656[63:48]     = Conv_out[165];
    assign  image_1_656[47:32]     = Conv_out[137];
    assign  image_1_656[31:16]     = Conv_out[136];
    assign  image_1_656[15:0]      = Conv_out[135];

    assign  image_1_657[143:128]   = Conv_out[196];
    assign  image_1_657[127:112]   = Conv_out[195];
    assign  image_1_657[111:96]    = Conv_out[194];
    assign  image_1_657[95:80]     = Conv_out[166];
    assign  image_1_657[79:64]     = Conv_out[165];
    assign  image_1_657[63:48]     = Conv_out[164];
    assign  image_1_657[47:32]     = Conv_out[136];
    assign  image_1_657[31:16]     = Conv_out[135];
    assign  image_1_657[15:0]      = Conv_out[134];

    assign  image_1_658[143:128]   = Conv_out[195];
    assign  image_1_658[127:112]   = Conv_out[194];
    assign  image_1_658[111:96]    = Conv_out[193];
    assign  image_1_658[95:80]     = Conv_out[165];
    assign  image_1_658[79:64]     = Conv_out[164];
    assign  image_1_658[63:48]     = Conv_out[163];
    assign  image_1_658[47:32]     = Conv_out[135];
    assign  image_1_658[31:16]     = Conv_out[134];
    assign  image_1_658[15:0]      = Conv_out[133];

    assign  image_1_659[143:128]   = Conv_out[194];
    assign  image_1_659[127:112]   = Conv_out[193];
    assign  image_1_659[111:96]    = Conv_out[192];
    assign  image_1_659[95:80]     = Conv_out[164];
    assign  image_1_659[79:64]     = Conv_out[163];
    assign  image_1_659[63:48]     = Conv_out[162];
    assign  image_1_659[47:32]     = Conv_out[134];
    assign  image_1_659[31:16]     = Conv_out[133];
    assign  image_1_659[15:0]      = Conv_out[132];

    assign  image_1_660[143:128]   = Conv_out[193];
    assign  image_1_660[127:112]   = Conv_out[192];
    assign  image_1_660[111:96]    = Conv_out[191];
    assign  image_1_660[95:80]     = Conv_out[163];
    assign  image_1_660[79:64]     = Conv_out[162];
    assign  image_1_660[63:48]     = Conv_out[161];
    assign  image_1_660[47:32]     = Conv_out[133];
    assign  image_1_660[31:16]     = Conv_out[132];
    assign  image_1_660[15:0]      = Conv_out[131];

    assign  image_1_661[143:128]   = Conv_out[192];
    assign  image_1_661[127:112]   = Conv_out[191];
    assign  image_1_661[111:96]    = Conv_out[190];
    assign  image_1_661[95:80]     = Conv_out[162];
    assign  image_1_661[79:64]     = Conv_out[161];
    assign  image_1_661[63:48]     = Conv_out[160];
    assign  image_1_661[47:32]     = Conv_out[132];
    assign  image_1_661[31:16]     = Conv_out[131];
    assign  image_1_661[15:0]      = Conv_out[130];

    assign  image_1_662[143:128]   = Conv_out[191];
    assign  image_1_662[127:112]   = Conv_out[190];
    assign  image_1_662[111:96]    = Conv_out[189];
    assign  image_1_662[95:80]     = Conv_out[161];
    assign  image_1_662[79:64]     = Conv_out[160];
    assign  image_1_662[63:48]     = Conv_out[159];
    assign  image_1_662[47:32]     = Conv_out[131];
    assign  image_1_662[31:16]     = Conv_out[130];
    assign  image_1_662[15:0]      = Conv_out[129];

    assign  image_1_663[143:128]   = Conv_out[190];
    assign  image_1_663[127:112]   = Conv_out[189];
    assign  image_1_663[111:96]    = Conv_out[188];
    assign  image_1_663[95:80]     = Conv_out[160];
    assign  image_1_663[79:64]     = Conv_out[159];
    assign  image_1_663[63:48]     = Conv_out[158];
    assign  image_1_663[47:32]     = Conv_out[130];
    assign  image_1_663[31:16]     = Conv_out[129];
    assign  image_1_663[15:0]      = Conv_out[128];

    assign  image_1_664[143:128]   = Conv_out[189];
    assign  image_1_664[127:112]   = Conv_out[188];
    assign  image_1_664[111:96]    = Conv_out[187];
    assign  image_1_664[95:80]     = Conv_out[159];
    assign  image_1_664[79:64]     = Conv_out[158];
    assign  image_1_664[63:48]     = Conv_out[157];
    assign  image_1_664[47:32]     = Conv_out[129];
    assign  image_1_664[31:16]     = Conv_out[128];
    assign  image_1_664[15:0]      = Conv_out[127];

    assign  image_1_665[143:128]   = Conv_out[188];
    assign  image_1_665[127:112]   = Conv_out[187];
    assign  image_1_665[111:96]    = Conv_out[186];
    assign  image_1_665[95:80]     = Conv_out[158];
    assign  image_1_665[79:64]     = Conv_out[157];
    assign  image_1_665[63:48]     = Conv_out[156];
    assign  image_1_665[47:32]     = Conv_out[128];
    assign  image_1_665[31:16]     = Conv_out[127];
    assign  image_1_665[15:0]      = Conv_out[126];

    assign  image_1_666[143:128]   = Conv_out[187];
    assign  image_1_666[127:112]   = Conv_out[186];
    assign  image_1_666[111:96]    = Conv_out[185];
    assign  image_1_666[95:80]     = Conv_out[157];
    assign  image_1_666[79:64]     = Conv_out[156];
    assign  image_1_666[63:48]     = Conv_out[155];
    assign  image_1_666[47:32]     = Conv_out[127];
    assign  image_1_666[31:16]     = Conv_out[126];
    assign  image_1_666[15:0]      = Conv_out[125];

    assign  image_1_667[143:128]   = Conv_out[186];
    assign  image_1_667[127:112]   = Conv_out[185];
    assign  image_1_667[111:96]    = Conv_out[184];
    assign  image_1_667[95:80]     = Conv_out[156];
    assign  image_1_667[79:64]     = Conv_out[155];
    assign  image_1_667[63:48]     = Conv_out[154];
    assign  image_1_667[47:32]     = Conv_out[126];
    assign  image_1_667[31:16]     = Conv_out[125];
    assign  image_1_667[15:0]      = Conv_out[124];

    assign  image_1_668[143:128]   = Conv_out[185];
    assign  image_1_668[127:112]   = Conv_out[184];
    assign  image_1_668[111:96]    = Conv_out[183];
    assign  image_1_668[95:80]     = Conv_out[155];
    assign  image_1_668[79:64]     = Conv_out[154];
    assign  image_1_668[63:48]     = Conv_out[153];
    assign  image_1_668[47:32]     = Conv_out[125];
    assign  image_1_668[31:16]     = Conv_out[124];
    assign  image_1_668[15:0]      = Conv_out[123];

    assign  image_1_669[143:128]   = Conv_out[184];
    assign  image_1_669[127:112]   = Conv_out[183];
    assign  image_1_669[111:96]    = Conv_out[182];
    assign  image_1_669[95:80]     = Conv_out[154];
    assign  image_1_669[79:64]     = Conv_out[153];
    assign  image_1_669[63:48]     = Conv_out[152];
    assign  image_1_669[47:32]     = Conv_out[124];
    assign  image_1_669[31:16]     = Conv_out[123];
    assign  image_1_669[15:0]      = Conv_out[122];

    assign  image_1_670[143:128]   = Conv_out[183];
    assign  image_1_670[127:112]   = Conv_out[182];
    assign  image_1_670[111:96]    = Conv_out[181];
    assign  image_1_670[95:80]     = Conv_out[153];
    assign  image_1_670[79:64]     = Conv_out[152];
    assign  image_1_670[63:48]     = Conv_out[151];
    assign  image_1_670[47:32]     = Conv_out[123];
    assign  image_1_670[31:16]     = Conv_out[122];
    assign  image_1_670[15:0]      = Conv_out[121];

    assign  image_1_671[143:128]   = Conv_out[182];
    assign  image_1_671[127:112]   = Conv_out[181];
    assign  image_1_671[111:96]    = Conv_out[180];
    assign  image_1_671[95:80]     = Conv_out[152];
    assign  image_1_671[79:64]     = Conv_out[151];
    assign  image_1_671[63:48]     = Conv_out[150];
    assign  image_1_671[47:32]     = Conv_out[122];
    assign  image_1_671[31:16]     = Conv_out[121];
    assign  image_1_671[15:0]      = Conv_out[120];

    assign  image_1_672[143:128]   = Conv_out[179];
    assign  image_1_672[127:112]   = Conv_out[178];
    assign  image_1_672[111:96]    = Conv_out[177];
    assign  image_1_672[95:80]     = Conv_out[149];
    assign  image_1_672[79:64]     = Conv_out[148];
    assign  image_1_672[63:48]     = Conv_out[147];
    assign  image_1_672[47:32]     = Conv_out[119];
    assign  image_1_672[31:16]     = Conv_out[118];
    assign  image_1_672[15:0]      = Conv_out[117];

    assign  image_1_673[143:128]   = Conv_out[178];
    assign  image_1_673[127:112]   = Conv_out[177];
    assign  image_1_673[111:96]    = Conv_out[176];
    assign  image_1_673[95:80]     = Conv_out[148];
    assign  image_1_673[79:64]     = Conv_out[147];
    assign  image_1_673[63:48]     = Conv_out[146];
    assign  image_1_673[47:32]     = Conv_out[118];
    assign  image_1_673[31:16]     = Conv_out[117];
    assign  image_1_673[15:0]      = Conv_out[116];

    assign  image_1_674[143:128]   = Conv_out[177];
    assign  image_1_674[127:112]   = Conv_out[176];
    assign  image_1_674[111:96]    = Conv_out[175];
    assign  image_1_674[95:80]     = Conv_out[147];
    assign  image_1_674[79:64]     = Conv_out[146];
    assign  image_1_674[63:48]     = Conv_out[145];
    assign  image_1_674[47:32]     = Conv_out[117];
    assign  image_1_674[31:16]     = Conv_out[116];
    assign  image_1_674[15:0]      = Conv_out[115];

    assign  image_1_675[143:128]   = Conv_out[176];
    assign  image_1_675[127:112]   = Conv_out[175];
    assign  image_1_675[111:96]    = Conv_out[174];
    assign  image_1_675[95:80]     = Conv_out[146];
    assign  image_1_675[79:64]     = Conv_out[145];
    assign  image_1_675[63:48]     = Conv_out[144];
    assign  image_1_675[47:32]     = Conv_out[116];
    assign  image_1_675[31:16]     = Conv_out[115];
    assign  image_1_675[15:0]      = Conv_out[114];

    assign  image_1_676[143:128]   = Conv_out[175];
    assign  image_1_676[127:112]   = Conv_out[174];
    assign  image_1_676[111:96]    = Conv_out[173];
    assign  image_1_676[95:80]     = Conv_out[145];
    assign  image_1_676[79:64]     = Conv_out[144];
    assign  image_1_676[63:48]     = Conv_out[143];
    assign  image_1_676[47:32]     = Conv_out[115];
    assign  image_1_676[31:16]     = Conv_out[114];
    assign  image_1_676[15:0]      = Conv_out[113];

    assign  image_1_677[143:128]   = Conv_out[174];
    assign  image_1_677[127:112]   = Conv_out[173];
    assign  image_1_677[111:96]    = Conv_out[172];
    assign  image_1_677[95:80]     = Conv_out[144];
    assign  image_1_677[79:64]     = Conv_out[143];
    assign  image_1_677[63:48]     = Conv_out[142];
    assign  image_1_677[47:32]     = Conv_out[114];
    assign  image_1_677[31:16]     = Conv_out[113];
    assign  image_1_677[15:0]      = Conv_out[112];

    assign  image_1_678[143:128]   = Conv_out[173];
    assign  image_1_678[127:112]   = Conv_out[172];
    assign  image_1_678[111:96]    = Conv_out[171];
    assign  image_1_678[95:80]     = Conv_out[143];
    assign  image_1_678[79:64]     = Conv_out[142];
    assign  image_1_678[63:48]     = Conv_out[141];
    assign  image_1_678[47:32]     = Conv_out[113];
    assign  image_1_678[31:16]     = Conv_out[112];
    assign  image_1_678[15:0]      = Conv_out[111];

    assign  image_1_679[143:128]   = Conv_out[172];
    assign  image_1_679[127:112]   = Conv_out[171];
    assign  image_1_679[111:96]    = Conv_out[170];
    assign  image_1_679[95:80]     = Conv_out[142];
    assign  image_1_679[79:64]     = Conv_out[141];
    assign  image_1_679[63:48]     = Conv_out[140];
    assign  image_1_679[47:32]     = Conv_out[112];
    assign  image_1_679[31:16]     = Conv_out[111];
    assign  image_1_679[15:0]      = Conv_out[110];

    assign  image_1_680[143:128]   = Conv_out[171];
    assign  image_1_680[127:112]   = Conv_out[170];
    assign  image_1_680[111:96]    = Conv_out[169];
    assign  image_1_680[95:80]     = Conv_out[141];
    assign  image_1_680[79:64]     = Conv_out[140];
    assign  image_1_680[63:48]     = Conv_out[139];
    assign  image_1_680[47:32]     = Conv_out[111];
    assign  image_1_680[31:16]     = Conv_out[110];
    assign  image_1_680[15:0]      = Conv_out[109];

    assign  image_1_681[143:128]   = Conv_out[170];
    assign  image_1_681[127:112]   = Conv_out[169];
    assign  image_1_681[111:96]    = Conv_out[168];
    assign  image_1_681[95:80]     = Conv_out[140];
    assign  image_1_681[79:64]     = Conv_out[139];
    assign  image_1_681[63:48]     = Conv_out[138];
    assign  image_1_681[47:32]     = Conv_out[110];
    assign  image_1_681[31:16]     = Conv_out[109];
    assign  image_1_681[15:0]      = Conv_out[108];

    assign  image_1_682[143:128]   = Conv_out[169];
    assign  image_1_682[127:112]   = Conv_out[168];
    assign  image_1_682[111:96]    = Conv_out[167];
    assign  image_1_682[95:80]     = Conv_out[139];
    assign  image_1_682[79:64]     = Conv_out[138];
    assign  image_1_682[63:48]     = Conv_out[137];
    assign  image_1_682[47:32]     = Conv_out[109];
    assign  image_1_682[31:16]     = Conv_out[108];
    assign  image_1_682[15:0]      = Conv_out[107];

    assign  image_1_683[143:128]   = Conv_out[168];
    assign  image_1_683[127:112]   = Conv_out[167];
    assign  image_1_683[111:96]    = Conv_out[166];
    assign  image_1_683[95:80]     = Conv_out[138];
    assign  image_1_683[79:64]     = Conv_out[137];
    assign  image_1_683[63:48]     = Conv_out[136];
    assign  image_1_683[47:32]     = Conv_out[108];
    assign  image_1_683[31:16]     = Conv_out[107];
    assign  image_1_683[15:0]      = Conv_out[106];

    assign  image_1_684[143:128]   = Conv_out[167];
    assign  image_1_684[127:112]   = Conv_out[166];
    assign  image_1_684[111:96]    = Conv_out[165];
    assign  image_1_684[95:80]     = Conv_out[137];
    assign  image_1_684[79:64]     = Conv_out[136];
    assign  image_1_684[63:48]     = Conv_out[135];
    assign  image_1_684[47:32]     = Conv_out[107];
    assign  image_1_684[31:16]     = Conv_out[106];
    assign  image_1_684[15:0]      = Conv_out[105];

    assign  image_1_685[143:128]   = Conv_out[166];
    assign  image_1_685[127:112]   = Conv_out[165];
    assign  image_1_685[111:96]    = Conv_out[164];
    assign  image_1_685[95:80]     = Conv_out[136];
    assign  image_1_685[79:64]     = Conv_out[135];
    assign  image_1_685[63:48]     = Conv_out[134];
    assign  image_1_685[47:32]     = Conv_out[106];
    assign  image_1_685[31:16]     = Conv_out[105];
    assign  image_1_685[15:0]      = Conv_out[104];

    assign  image_1_686[143:128]   = Conv_out[165];
    assign  image_1_686[127:112]   = Conv_out[164];
    assign  image_1_686[111:96]    = Conv_out[163];
    assign  image_1_686[95:80]     = Conv_out[135];
    assign  image_1_686[79:64]     = Conv_out[134];
    assign  image_1_686[63:48]     = Conv_out[133];
    assign  image_1_686[47:32]     = Conv_out[105];
    assign  image_1_686[31:16]     = Conv_out[104];
    assign  image_1_686[15:0]      = Conv_out[103];

    assign  image_1_687[143:128]   = Conv_out[164];
    assign  image_1_687[127:112]   = Conv_out[163];
    assign  image_1_687[111:96]    = Conv_out[162];
    assign  image_1_687[95:80]     = Conv_out[134];
    assign  image_1_687[79:64]     = Conv_out[133];
    assign  image_1_687[63:48]     = Conv_out[132];
    assign  image_1_687[47:32]     = Conv_out[104];
    assign  image_1_687[31:16]     = Conv_out[103];
    assign  image_1_687[15:0]      = Conv_out[102];

    assign  image_1_688[143:128]   = Conv_out[163];
    assign  image_1_688[127:112]   = Conv_out[162];
    assign  image_1_688[111:96]    = Conv_out[161];
    assign  image_1_688[95:80]     = Conv_out[133];
    assign  image_1_688[79:64]     = Conv_out[132];
    assign  image_1_688[63:48]     = Conv_out[131];
    assign  image_1_688[47:32]     = Conv_out[103];
    assign  image_1_688[31:16]     = Conv_out[102];
    assign  image_1_688[15:0]      = Conv_out[101];

    assign  image_1_689[143:128]   = Conv_out[162];
    assign  image_1_689[127:112]   = Conv_out[161];
    assign  image_1_689[111:96]    = Conv_out[160];
    assign  image_1_689[95:80]     = Conv_out[132];
    assign  image_1_689[79:64]     = Conv_out[131];
    assign  image_1_689[63:48]     = Conv_out[130];
    assign  image_1_689[47:32]     = Conv_out[102];
    assign  image_1_689[31:16]     = Conv_out[101];
    assign  image_1_689[15:0]      = Conv_out[100];

    assign  image_1_690[143:128]   = Conv_out[161];
    assign  image_1_690[127:112]   = Conv_out[160];
    assign  image_1_690[111:96]    = Conv_out[159];
    assign  image_1_690[95:80]     = Conv_out[131];
    assign  image_1_690[79:64]     = Conv_out[130];
    assign  image_1_690[63:48]     = Conv_out[129];
    assign  image_1_690[47:32]     = Conv_out[101];
    assign  image_1_690[31:16]     = Conv_out[100];
    assign  image_1_690[15:0]      = Conv_out[99];

    assign  image_1_691[143:128]   = Conv_out[160];
    assign  image_1_691[127:112]   = Conv_out[159];
    assign  image_1_691[111:96]    = Conv_out[158];
    assign  image_1_691[95:80]     = Conv_out[130];
    assign  image_1_691[79:64]     = Conv_out[129];
    assign  image_1_691[63:48]     = Conv_out[128];
    assign  image_1_691[47:32]     = Conv_out[100];
    assign  image_1_691[31:16]     = Conv_out[99];
    assign  image_1_691[15:0]      = Conv_out[98];

    assign  image_1_692[143:128]   = Conv_out[159];
    assign  image_1_692[127:112]   = Conv_out[158];
    assign  image_1_692[111:96]    = Conv_out[157];
    assign  image_1_692[95:80]     = Conv_out[129];
    assign  image_1_692[79:64]     = Conv_out[128];
    assign  image_1_692[63:48]     = Conv_out[127];
    assign  image_1_692[47:32]     = Conv_out[99];
    assign  image_1_692[31:16]     = Conv_out[98];
    assign  image_1_692[15:0]      = Conv_out[97];

    assign  image_1_693[143:128]   = Conv_out[158];
    assign  image_1_693[127:112]   = Conv_out[157];
    assign  image_1_693[111:96]    = Conv_out[156];
    assign  image_1_693[95:80]     = Conv_out[128];
    assign  image_1_693[79:64]     = Conv_out[127];
    assign  image_1_693[63:48]     = Conv_out[126];
    assign  image_1_693[47:32]     = Conv_out[98];
    assign  image_1_693[31:16]     = Conv_out[97];
    assign  image_1_693[15:0]      = Conv_out[96];

    assign  image_1_694[143:128]   = Conv_out[157];
    assign  image_1_694[127:112]   = Conv_out[156];
    assign  image_1_694[111:96]    = Conv_out[155];
    assign  image_1_694[95:80]     = Conv_out[127];
    assign  image_1_694[79:64]     = Conv_out[126];
    assign  image_1_694[63:48]     = Conv_out[125];
    assign  image_1_694[47:32]     = Conv_out[97];
    assign  image_1_694[31:16]     = Conv_out[96];
    assign  image_1_694[15:0]      = Conv_out[95];

    assign  image_1_695[143:128]   = Conv_out[156];
    assign  image_1_695[127:112]   = Conv_out[155];
    assign  image_1_695[111:96]    = Conv_out[154];
    assign  image_1_695[95:80]     = Conv_out[126];
    assign  image_1_695[79:64]     = Conv_out[125];
    assign  image_1_695[63:48]     = Conv_out[124];
    assign  image_1_695[47:32]     = Conv_out[96];
    assign  image_1_695[31:16]     = Conv_out[95];
    assign  image_1_695[15:0]      = Conv_out[94];

    assign  image_1_696[143:128]   = Conv_out[155];
    assign  image_1_696[127:112]   = Conv_out[154];
    assign  image_1_696[111:96]    = Conv_out[153];
    assign  image_1_696[95:80]     = Conv_out[125];
    assign  image_1_696[79:64]     = Conv_out[124];
    assign  image_1_696[63:48]     = Conv_out[123];
    assign  image_1_696[47:32]     = Conv_out[95];
    assign  image_1_696[31:16]     = Conv_out[94];
    assign  image_1_696[15:0]      = Conv_out[93];

    assign  image_1_697[143:128]   = Conv_out[154];
    assign  image_1_697[127:112]   = Conv_out[153];
    assign  image_1_697[111:96]    = Conv_out[152];
    assign  image_1_697[95:80]     = Conv_out[124];
    assign  image_1_697[79:64]     = Conv_out[123];
    assign  image_1_697[63:48]     = Conv_out[122];
    assign  image_1_697[47:32]     = Conv_out[94];
    assign  image_1_697[31:16]     = Conv_out[93];
    assign  image_1_697[15:0]      = Conv_out[92];

    assign  image_1_698[143:128]   = Conv_out[153];
    assign  image_1_698[127:112]   = Conv_out[152];
    assign  image_1_698[111:96]    = Conv_out[151];
    assign  image_1_698[95:80]     = Conv_out[123];
    assign  image_1_698[79:64]     = Conv_out[122];
    assign  image_1_698[63:48]     = Conv_out[121];
    assign  image_1_698[47:32]     = Conv_out[93];
    assign  image_1_698[31:16]     = Conv_out[92];
    assign  image_1_698[15:0]      = Conv_out[91];

    assign  image_1_699[143:128]   = Conv_out[152];
    assign  image_1_699[127:112]   = Conv_out[151];
    assign  image_1_699[111:96]    = Conv_out[150];
    assign  image_1_699[95:80]     = Conv_out[122];
    assign  image_1_699[79:64]     = Conv_out[121];
    assign  image_1_699[63:48]     = Conv_out[120];
    assign  image_1_699[47:32]     = Conv_out[92];
    assign  image_1_699[31:16]     = Conv_out[91];
    assign  image_1_699[15:0]      = Conv_out[90];

    assign  image_1_700[143:128]   = Conv_out[149];
    assign  image_1_700[127:112]   = Conv_out[148];
    assign  image_1_700[111:96]    = Conv_out[147];
    assign  image_1_700[95:80]     = Conv_out[119];
    assign  image_1_700[79:64]     = Conv_out[118];
    assign  image_1_700[63:48]     = Conv_out[117];
    assign  image_1_700[47:32]     = Conv_out[89];
    assign  image_1_700[31:16]     = Conv_out[88];
    assign  image_1_700[15:0]      = Conv_out[87];

    assign  image_1_701[143:128]   = Conv_out[148];
    assign  image_1_701[127:112]   = Conv_out[147];
    assign  image_1_701[111:96]    = Conv_out[146];
    assign  image_1_701[95:80]     = Conv_out[118];
    assign  image_1_701[79:64]     = Conv_out[117];
    assign  image_1_701[63:48]     = Conv_out[116];
    assign  image_1_701[47:32]     = Conv_out[88];
    assign  image_1_701[31:16]     = Conv_out[87];
    assign  image_1_701[15:0]      = Conv_out[86];

    assign  image_1_702[143:128]   = Conv_out[147];
    assign  image_1_702[127:112]   = Conv_out[146];
    assign  image_1_702[111:96]    = Conv_out[145];
    assign  image_1_702[95:80]     = Conv_out[117];
    assign  image_1_702[79:64]     = Conv_out[116];
    assign  image_1_702[63:48]     = Conv_out[115];
    assign  image_1_702[47:32]     = Conv_out[87];
    assign  image_1_702[31:16]     = Conv_out[86];
    assign  image_1_702[15:0]      = Conv_out[85];

    assign  image_1_703[143:128]   = Conv_out[146];
    assign  image_1_703[127:112]   = Conv_out[145];
    assign  image_1_703[111:96]    = Conv_out[144];
    assign  image_1_703[95:80]     = Conv_out[116];
    assign  image_1_703[79:64]     = Conv_out[115];
    assign  image_1_703[63:48]     = Conv_out[114];
    assign  image_1_703[47:32]     = Conv_out[86];
    assign  image_1_703[31:16]     = Conv_out[85];
    assign  image_1_703[15:0]      = Conv_out[84];

    assign  image_1_704[143:128]   = Conv_out[145];
    assign  image_1_704[127:112]   = Conv_out[144];
    assign  image_1_704[111:96]    = Conv_out[143];
    assign  image_1_704[95:80]     = Conv_out[115];
    assign  image_1_704[79:64]     = Conv_out[114];
    assign  image_1_704[63:48]     = Conv_out[113];
    assign  image_1_704[47:32]     = Conv_out[85];
    assign  image_1_704[31:16]     = Conv_out[84];
    assign  image_1_704[15:0]      = Conv_out[83];

    assign  image_1_705[143:128]   = Conv_out[144];
    assign  image_1_705[127:112]   = Conv_out[143];
    assign  image_1_705[111:96]    = Conv_out[142];
    assign  image_1_705[95:80]     = Conv_out[114];
    assign  image_1_705[79:64]     = Conv_out[113];
    assign  image_1_705[63:48]     = Conv_out[112];
    assign  image_1_705[47:32]     = Conv_out[84];
    assign  image_1_705[31:16]     = Conv_out[83];
    assign  image_1_705[15:0]      = Conv_out[82];

    assign  image_1_706[143:128]   = Conv_out[143];
    assign  image_1_706[127:112]   = Conv_out[142];
    assign  image_1_706[111:96]    = Conv_out[141];
    assign  image_1_706[95:80]     = Conv_out[113];
    assign  image_1_706[79:64]     = Conv_out[112];
    assign  image_1_706[63:48]     = Conv_out[111];
    assign  image_1_706[47:32]     = Conv_out[83];
    assign  image_1_706[31:16]     = Conv_out[82];
    assign  image_1_706[15:0]      = Conv_out[81];

    assign  image_1_707[143:128]   = Conv_out[142];
    assign  image_1_707[127:112]   = Conv_out[141];
    assign  image_1_707[111:96]    = Conv_out[140];
    assign  image_1_707[95:80]     = Conv_out[112];
    assign  image_1_707[79:64]     = Conv_out[111];
    assign  image_1_707[63:48]     = Conv_out[110];
    assign  image_1_707[47:32]     = Conv_out[82];
    assign  image_1_707[31:16]     = Conv_out[81];
    assign  image_1_707[15:0]      = Conv_out[80];

    assign  image_1_708[143:128]   = Conv_out[141];
    assign  image_1_708[127:112]   = Conv_out[140];
    assign  image_1_708[111:96]    = Conv_out[139];
    assign  image_1_708[95:80]     = Conv_out[111];
    assign  image_1_708[79:64]     = Conv_out[110];
    assign  image_1_708[63:48]     = Conv_out[109];
    assign  image_1_708[47:32]     = Conv_out[81];
    assign  image_1_708[31:16]     = Conv_out[80];
    assign  image_1_708[15:0]      = Conv_out[79];

    assign  image_1_709[143:128]   = Conv_out[140];
    assign  image_1_709[127:112]   = Conv_out[139];
    assign  image_1_709[111:96]    = Conv_out[138];
    assign  image_1_709[95:80]     = Conv_out[110];
    assign  image_1_709[79:64]     = Conv_out[109];
    assign  image_1_709[63:48]     = Conv_out[108];
    assign  image_1_709[47:32]     = Conv_out[80];
    assign  image_1_709[31:16]     = Conv_out[79];
    assign  image_1_709[15:0]      = Conv_out[78];

    assign  image_1_710[143:128]   = Conv_out[139];
    assign  image_1_710[127:112]   = Conv_out[138];
    assign  image_1_710[111:96]    = Conv_out[137];
    assign  image_1_710[95:80]     = Conv_out[109];
    assign  image_1_710[79:64]     = Conv_out[108];
    assign  image_1_710[63:48]     = Conv_out[107];
    assign  image_1_710[47:32]     = Conv_out[79];
    assign  image_1_710[31:16]     = Conv_out[78];
    assign  image_1_710[15:0]      = Conv_out[77];

    assign  image_1_711[143:128]   = Conv_out[138];
    assign  image_1_711[127:112]   = Conv_out[137];
    assign  image_1_711[111:96]    = Conv_out[136];
    assign  image_1_711[95:80]     = Conv_out[108];
    assign  image_1_711[79:64]     = Conv_out[107];
    assign  image_1_711[63:48]     = Conv_out[106];
    assign  image_1_711[47:32]     = Conv_out[78];
    assign  image_1_711[31:16]     = Conv_out[77];
    assign  image_1_711[15:0]      = Conv_out[76];

    assign  image_1_712[143:128]   = Conv_out[137];
    assign  image_1_712[127:112]   = Conv_out[136];
    assign  image_1_712[111:96]    = Conv_out[135];
    assign  image_1_712[95:80]     = Conv_out[107];
    assign  image_1_712[79:64]     = Conv_out[106];
    assign  image_1_712[63:48]     = Conv_out[105];
    assign  image_1_712[47:32]     = Conv_out[77];
    assign  image_1_712[31:16]     = Conv_out[76];
    assign  image_1_712[15:0]      = Conv_out[75];

    assign  image_1_713[143:128]   = Conv_out[136];
    assign  image_1_713[127:112]   = Conv_out[135];
    assign  image_1_713[111:96]    = Conv_out[134];
    assign  image_1_713[95:80]     = Conv_out[106];
    assign  image_1_713[79:64]     = Conv_out[105];
    assign  image_1_713[63:48]     = Conv_out[104];
    assign  image_1_713[47:32]     = Conv_out[76];
    assign  image_1_713[31:16]     = Conv_out[75];
    assign  image_1_713[15:0]      = Conv_out[74];

    assign  image_1_714[143:128]   = Conv_out[135];
    assign  image_1_714[127:112]   = Conv_out[134];
    assign  image_1_714[111:96]    = Conv_out[133];
    assign  image_1_714[95:80]     = Conv_out[105];
    assign  image_1_714[79:64]     = Conv_out[104];
    assign  image_1_714[63:48]     = Conv_out[103];
    assign  image_1_714[47:32]     = Conv_out[75];
    assign  image_1_714[31:16]     = Conv_out[74];
    assign  image_1_714[15:0]      = Conv_out[73];

    assign  image_1_715[143:128]   = Conv_out[134];
    assign  image_1_715[127:112]   = Conv_out[133];
    assign  image_1_715[111:96]    = Conv_out[132];
    assign  image_1_715[95:80]     = Conv_out[104];
    assign  image_1_715[79:64]     = Conv_out[103];
    assign  image_1_715[63:48]     = Conv_out[102];
    assign  image_1_715[47:32]     = Conv_out[74];
    assign  image_1_715[31:16]     = Conv_out[73];
    assign  image_1_715[15:0]      = Conv_out[72];

    assign  image_1_716[143:128]   = Conv_out[133];
    assign  image_1_716[127:112]   = Conv_out[132];
    assign  image_1_716[111:96]    = Conv_out[131];
    assign  image_1_716[95:80]     = Conv_out[103];
    assign  image_1_716[79:64]     = Conv_out[102];
    assign  image_1_716[63:48]     = Conv_out[101];
    assign  image_1_716[47:32]     = Conv_out[73];
    assign  image_1_716[31:16]     = Conv_out[72];
    assign  image_1_716[15:0]      = Conv_out[71];

    assign  image_1_717[143:128]   = Conv_out[132];
    assign  image_1_717[127:112]   = Conv_out[131];
    assign  image_1_717[111:96]    = Conv_out[130];
    assign  image_1_717[95:80]     = Conv_out[102];
    assign  image_1_717[79:64]     = Conv_out[101];
    assign  image_1_717[63:48]     = Conv_out[100];
    assign  image_1_717[47:32]     = Conv_out[72];
    assign  image_1_717[31:16]     = Conv_out[71];
    assign  image_1_717[15:0]      = Conv_out[70];

    assign  image_1_718[143:128]   = Conv_out[131];
    assign  image_1_718[127:112]   = Conv_out[130];
    assign  image_1_718[111:96]    = Conv_out[129];
    assign  image_1_718[95:80]     = Conv_out[101];
    assign  image_1_718[79:64]     = Conv_out[100];
    assign  image_1_718[63:48]     = Conv_out[99];
    assign  image_1_718[47:32]     = Conv_out[71];
    assign  image_1_718[31:16]     = Conv_out[70];
    assign  image_1_718[15:0]      = Conv_out[69];

    assign  image_1_719[143:128]   = Conv_out[130];
    assign  image_1_719[127:112]   = Conv_out[129];
    assign  image_1_719[111:96]    = Conv_out[128];
    assign  image_1_719[95:80]     = Conv_out[100];
    assign  image_1_719[79:64]     = Conv_out[99];
    assign  image_1_719[63:48]     = Conv_out[98];
    assign  image_1_719[47:32]     = Conv_out[70];
    assign  image_1_719[31:16]     = Conv_out[69];
    assign  image_1_719[15:0]      = Conv_out[68];

    assign  image_1_720[143:128]   = Conv_out[129];
    assign  image_1_720[127:112]   = Conv_out[128];
    assign  image_1_720[111:96]    = Conv_out[127];
    assign  image_1_720[95:80]     = Conv_out[99];
    assign  image_1_720[79:64]     = Conv_out[98];
    assign  image_1_720[63:48]     = Conv_out[97];
    assign  image_1_720[47:32]     = Conv_out[69];
    assign  image_1_720[31:16]     = Conv_out[68];
    assign  image_1_720[15:0]      = Conv_out[67];

    assign  image_1_721[143:128]   = Conv_out[128];
    assign  image_1_721[127:112]   = Conv_out[127];
    assign  image_1_721[111:96]    = Conv_out[126];
    assign  image_1_721[95:80]     = Conv_out[98];
    assign  image_1_721[79:64]     = Conv_out[97];
    assign  image_1_721[63:48]     = Conv_out[96];
    assign  image_1_721[47:32]     = Conv_out[68];
    assign  image_1_721[31:16]     = Conv_out[67];
    assign  image_1_721[15:0]      = Conv_out[66];

    assign  image_1_722[143:128]   = Conv_out[127];
    assign  image_1_722[127:112]   = Conv_out[126];
    assign  image_1_722[111:96]    = Conv_out[125];
    assign  image_1_722[95:80]     = Conv_out[97];
    assign  image_1_722[79:64]     = Conv_out[96];
    assign  image_1_722[63:48]     = Conv_out[95];
    assign  image_1_722[47:32]     = Conv_out[67];
    assign  image_1_722[31:16]     = Conv_out[66];
    assign  image_1_722[15:0]      = Conv_out[65];

    assign  image_1_723[143:128]   = Conv_out[126];
    assign  image_1_723[127:112]   = Conv_out[125];
    assign  image_1_723[111:96]    = Conv_out[124];
    assign  image_1_723[95:80]     = Conv_out[96];
    assign  image_1_723[79:64]     = Conv_out[95];
    assign  image_1_723[63:48]     = Conv_out[94];
    assign  image_1_723[47:32]     = Conv_out[66];
    assign  image_1_723[31:16]     = Conv_out[65];
    assign  image_1_723[15:0]      = Conv_out[64];

    assign  image_1_724[143:128]   = Conv_out[125];
    assign  image_1_724[127:112]   = Conv_out[124];
    assign  image_1_724[111:96]    = Conv_out[123];
    assign  image_1_724[95:80]     = Conv_out[95];
    assign  image_1_724[79:64]     = Conv_out[94];
    assign  image_1_724[63:48]     = Conv_out[93];
    assign  image_1_724[47:32]     = Conv_out[65];
    assign  image_1_724[31:16]     = Conv_out[64];
    assign  image_1_724[15:0]      = Conv_out[63];

    assign  image_1_725[143:128]   = Conv_out[124];
    assign  image_1_725[127:112]   = Conv_out[123];
    assign  image_1_725[111:96]    = Conv_out[122];
    assign  image_1_725[95:80]     = Conv_out[94];
    assign  image_1_725[79:64]     = Conv_out[93];
    assign  image_1_725[63:48]     = Conv_out[92];
    assign  image_1_725[47:32]     = Conv_out[64];
    assign  image_1_725[31:16]     = Conv_out[63];
    assign  image_1_725[15:0]      = Conv_out[62];

    assign  image_1_726[143:128]   = Conv_out[123];
    assign  image_1_726[127:112]   = Conv_out[122];
    assign  image_1_726[111:96]    = Conv_out[121];
    assign  image_1_726[95:80]     = Conv_out[93];
    assign  image_1_726[79:64]     = Conv_out[92];
    assign  image_1_726[63:48]     = Conv_out[91];
    assign  image_1_726[47:32]     = Conv_out[63];
    assign  image_1_726[31:16]     = Conv_out[62];
    assign  image_1_726[15:0]      = Conv_out[61];

    assign  image_1_727[143:128]   = Conv_out[122];
    assign  image_1_727[127:112]   = Conv_out[121];
    assign  image_1_727[111:96]    = Conv_out[120];
    assign  image_1_727[95:80]     = Conv_out[92];
    assign  image_1_727[79:64]     = Conv_out[91];
    assign  image_1_727[63:48]     = Conv_out[90];
    assign  image_1_727[47:32]     = Conv_out[62];
    assign  image_1_727[31:16]     = Conv_out[61];
    assign  image_1_727[15:0]      = Conv_out[60];

    assign  image_1_728[143:128]   = Conv_out[119];
    assign  image_1_728[127:112]   = Conv_out[118];
    assign  image_1_728[111:96]    = Conv_out[117];
    assign  image_1_728[95:80]     = Conv_out[89];
    assign  image_1_728[79:64]     = Conv_out[88];
    assign  image_1_728[63:48]     = Conv_out[87];
    assign  image_1_728[47:32]     = Conv_out[59];
    assign  image_1_728[31:16]     = Conv_out[58];
    assign  image_1_728[15:0]      = Conv_out[57];

    assign  image_1_729[143:128]   = Conv_out[118];
    assign  image_1_729[127:112]   = Conv_out[117];
    assign  image_1_729[111:96]    = Conv_out[116];
    assign  image_1_729[95:80]     = Conv_out[88];
    assign  image_1_729[79:64]     = Conv_out[87];
    assign  image_1_729[63:48]     = Conv_out[86];
    assign  image_1_729[47:32]     = Conv_out[58];
    assign  image_1_729[31:16]     = Conv_out[57];
    assign  image_1_729[15:0]      = Conv_out[56];

    assign  image_1_730[143:128]   = Conv_out[117];
    assign  image_1_730[127:112]   = Conv_out[116];
    assign  image_1_730[111:96]    = Conv_out[115];
    assign  image_1_730[95:80]     = Conv_out[87];
    assign  image_1_730[79:64]     = Conv_out[86];
    assign  image_1_730[63:48]     = Conv_out[85];
    assign  image_1_730[47:32]     = Conv_out[57];
    assign  image_1_730[31:16]     = Conv_out[56];
    assign  image_1_730[15:0]      = Conv_out[55];

    assign  image_1_731[143:128]   = Conv_out[116];
    assign  image_1_731[127:112]   = Conv_out[115];
    assign  image_1_731[111:96]    = Conv_out[114];
    assign  image_1_731[95:80]     = Conv_out[86];
    assign  image_1_731[79:64]     = Conv_out[85];
    assign  image_1_731[63:48]     = Conv_out[84];
    assign  image_1_731[47:32]     = Conv_out[56];
    assign  image_1_731[31:16]     = Conv_out[55];
    assign  image_1_731[15:0]      = Conv_out[54];

    assign  image_1_732[143:128]   = Conv_out[115];
    assign  image_1_732[127:112]   = Conv_out[114];
    assign  image_1_732[111:96]    = Conv_out[113];
    assign  image_1_732[95:80]     = Conv_out[85];
    assign  image_1_732[79:64]     = Conv_out[84];
    assign  image_1_732[63:48]     = Conv_out[83];
    assign  image_1_732[47:32]     = Conv_out[55];
    assign  image_1_732[31:16]     = Conv_out[54];
    assign  image_1_732[15:0]      = Conv_out[53];

    assign  image_1_733[143:128]   = Conv_out[114];
    assign  image_1_733[127:112]   = Conv_out[113];
    assign  image_1_733[111:96]    = Conv_out[112];
    assign  image_1_733[95:80]     = Conv_out[84];
    assign  image_1_733[79:64]     = Conv_out[83];
    assign  image_1_733[63:48]     = Conv_out[82];
    assign  image_1_733[47:32]     = Conv_out[54];
    assign  image_1_733[31:16]     = Conv_out[53];
    assign  image_1_733[15:0]      = Conv_out[52];

    assign  image_1_734[143:128]   = Conv_out[113];
    assign  image_1_734[127:112]   = Conv_out[112];
    assign  image_1_734[111:96]    = Conv_out[111];
    assign  image_1_734[95:80]     = Conv_out[83];
    assign  image_1_734[79:64]     = Conv_out[82];
    assign  image_1_734[63:48]     = Conv_out[81];
    assign  image_1_734[47:32]     = Conv_out[53];
    assign  image_1_734[31:16]     = Conv_out[52];
    assign  image_1_734[15:0]      = Conv_out[51];

    assign  image_1_735[143:128]   = Conv_out[112];
    assign  image_1_735[127:112]   = Conv_out[111];
    assign  image_1_735[111:96]    = Conv_out[110];
    assign  image_1_735[95:80]     = Conv_out[82];
    assign  image_1_735[79:64]     = Conv_out[81];
    assign  image_1_735[63:48]     = Conv_out[80];
    assign  image_1_735[47:32]     = Conv_out[52];
    assign  image_1_735[31:16]     = Conv_out[51];
    assign  image_1_735[15:0]      = Conv_out[50];

    assign  image_1_736[143:128]   = Conv_out[111];
    assign  image_1_736[127:112]   = Conv_out[110];
    assign  image_1_736[111:96]    = Conv_out[109];
    assign  image_1_736[95:80]     = Conv_out[81];
    assign  image_1_736[79:64]     = Conv_out[80];
    assign  image_1_736[63:48]     = Conv_out[79];
    assign  image_1_736[47:32]     = Conv_out[51];
    assign  image_1_736[31:16]     = Conv_out[50];
    assign  image_1_736[15:0]      = Conv_out[49];

    assign  image_1_737[143:128]   = Conv_out[110];
    assign  image_1_737[127:112]   = Conv_out[109];
    assign  image_1_737[111:96]    = Conv_out[108];
    assign  image_1_737[95:80]     = Conv_out[80];
    assign  image_1_737[79:64]     = Conv_out[79];
    assign  image_1_737[63:48]     = Conv_out[78];
    assign  image_1_737[47:32]     = Conv_out[50];
    assign  image_1_737[31:16]     = Conv_out[49];
    assign  image_1_737[15:0]      = Conv_out[48];

    assign  image_1_738[143:128]   = Conv_out[109];
    assign  image_1_738[127:112]   = Conv_out[108];
    assign  image_1_738[111:96]    = Conv_out[107];
    assign  image_1_738[95:80]     = Conv_out[79];
    assign  image_1_738[79:64]     = Conv_out[78];
    assign  image_1_738[63:48]     = Conv_out[77];
    assign  image_1_738[47:32]     = Conv_out[49];
    assign  image_1_738[31:16]     = Conv_out[48];
    assign  image_1_738[15:0]      = Conv_out[47];

    assign  image_1_739[143:128]   = Conv_out[108];
    assign  image_1_739[127:112]   = Conv_out[107];
    assign  image_1_739[111:96]    = Conv_out[106];
    assign  image_1_739[95:80]     = Conv_out[78];
    assign  image_1_739[79:64]     = Conv_out[77];
    assign  image_1_739[63:48]     = Conv_out[76];
    assign  image_1_739[47:32]     = Conv_out[48];
    assign  image_1_739[31:16]     = Conv_out[47];
    assign  image_1_739[15:0]      = Conv_out[46];

    assign  image_1_740[143:128]   = Conv_out[107];
    assign  image_1_740[127:112]   = Conv_out[106];
    assign  image_1_740[111:96]    = Conv_out[105];
    assign  image_1_740[95:80]     = Conv_out[77];
    assign  image_1_740[79:64]     = Conv_out[76];
    assign  image_1_740[63:48]     = Conv_out[75];
    assign  image_1_740[47:32]     = Conv_out[47];
    assign  image_1_740[31:16]     = Conv_out[46];
    assign  image_1_740[15:0]      = Conv_out[45];

    assign  image_1_741[143:128]   = Conv_out[106];
    assign  image_1_741[127:112]   = Conv_out[105];
    assign  image_1_741[111:96]    = Conv_out[104];
    assign  image_1_741[95:80]     = Conv_out[76];
    assign  image_1_741[79:64]     = Conv_out[75];
    assign  image_1_741[63:48]     = Conv_out[74];
    assign  image_1_741[47:32]     = Conv_out[46];
    assign  image_1_741[31:16]     = Conv_out[45];
    assign  image_1_741[15:0]      = Conv_out[44];

    assign  image_1_742[143:128]   = Conv_out[105];
    assign  image_1_742[127:112]   = Conv_out[104];
    assign  image_1_742[111:96]    = Conv_out[103];
    assign  image_1_742[95:80]     = Conv_out[75];
    assign  image_1_742[79:64]     = Conv_out[74];
    assign  image_1_742[63:48]     = Conv_out[73];
    assign  image_1_742[47:32]     = Conv_out[45];
    assign  image_1_742[31:16]     = Conv_out[44];
    assign  image_1_742[15:0]      = Conv_out[43];

    assign  image_1_743[143:128]   = Conv_out[104];
    assign  image_1_743[127:112]   = Conv_out[103];
    assign  image_1_743[111:96]    = Conv_out[102];
    assign  image_1_743[95:80]     = Conv_out[74];
    assign  image_1_743[79:64]     = Conv_out[73];
    assign  image_1_743[63:48]     = Conv_out[72];
    assign  image_1_743[47:32]     = Conv_out[44];
    assign  image_1_743[31:16]     = Conv_out[43];
    assign  image_1_743[15:0]      = Conv_out[42];

    assign  image_1_744[143:128]   = Conv_out[103];
    assign  image_1_744[127:112]   = Conv_out[102];
    assign  image_1_744[111:96]    = Conv_out[101];
    assign  image_1_744[95:80]     = Conv_out[73];
    assign  image_1_744[79:64]     = Conv_out[72];
    assign  image_1_744[63:48]     = Conv_out[71];
    assign  image_1_744[47:32]     = Conv_out[43];
    assign  image_1_744[31:16]     = Conv_out[42];
    assign  image_1_744[15:0]      = Conv_out[41];

    assign  image_1_745[143:128]   = Conv_out[102];
    assign  image_1_745[127:112]   = Conv_out[101];
    assign  image_1_745[111:96]    = Conv_out[100];
    assign  image_1_745[95:80]     = Conv_out[72];
    assign  image_1_745[79:64]     = Conv_out[71];
    assign  image_1_745[63:48]     = Conv_out[70];
    assign  image_1_745[47:32]     = Conv_out[42];
    assign  image_1_745[31:16]     = Conv_out[41];
    assign  image_1_745[15:0]      = Conv_out[40];

    assign  image_1_746[143:128]   = Conv_out[101];
    assign  image_1_746[127:112]   = Conv_out[100];
    assign  image_1_746[111:96]    = Conv_out[99];
    assign  image_1_746[95:80]     = Conv_out[71];
    assign  image_1_746[79:64]     = Conv_out[70];
    assign  image_1_746[63:48]     = Conv_out[69];
    assign  image_1_746[47:32]     = Conv_out[41];
    assign  image_1_746[31:16]     = Conv_out[40];
    assign  image_1_746[15:0]      = Conv_out[39];

    assign  image_1_747[143:128]   = Conv_out[100];
    assign  image_1_747[127:112]   = Conv_out[99];
    assign  image_1_747[111:96]    = Conv_out[98];
    assign  image_1_747[95:80]     = Conv_out[70];
    assign  image_1_747[79:64]     = Conv_out[69];
    assign  image_1_747[63:48]     = Conv_out[68];
    assign  image_1_747[47:32]     = Conv_out[40];
    assign  image_1_747[31:16]     = Conv_out[39];
    assign  image_1_747[15:0]      = Conv_out[38];

    assign  image_1_748[143:128]   = Conv_out[99];
    assign  image_1_748[127:112]   = Conv_out[98];
    assign  image_1_748[111:96]    = Conv_out[97];
    assign  image_1_748[95:80]     = Conv_out[69];
    assign  image_1_748[79:64]     = Conv_out[68];
    assign  image_1_748[63:48]     = Conv_out[67];
    assign  image_1_748[47:32]     = Conv_out[39];
    assign  image_1_748[31:16]     = Conv_out[38];
    assign  image_1_748[15:0]      = Conv_out[37];

    assign  image_1_749[143:128]   = Conv_out[98];
    assign  image_1_749[127:112]   = Conv_out[97];
    assign  image_1_749[111:96]    = Conv_out[96];
    assign  image_1_749[95:80]     = Conv_out[68];
    assign  image_1_749[79:64]     = Conv_out[67];
    assign  image_1_749[63:48]     = Conv_out[66];
    assign  image_1_749[47:32]     = Conv_out[38];
    assign  image_1_749[31:16]     = Conv_out[37];
    assign  image_1_749[15:0]      = Conv_out[36];

    assign  image_1_750[143:128]   = Conv_out[97];
    assign  image_1_750[127:112]   = Conv_out[96];
    assign  image_1_750[111:96]    = Conv_out[95];
    assign  image_1_750[95:80]     = Conv_out[67];
    assign  image_1_750[79:64]     = Conv_out[66];
    assign  image_1_750[63:48]     = Conv_out[65];
    assign  image_1_750[47:32]     = Conv_out[37];
    assign  image_1_750[31:16]     = Conv_out[36];
    assign  image_1_750[15:0]      = Conv_out[35];

    assign  image_1_751[143:128]   = Conv_out[96];
    assign  image_1_751[127:112]   = Conv_out[95];
    assign  image_1_751[111:96]    = Conv_out[94];
    assign  image_1_751[95:80]     = Conv_out[66];
    assign  image_1_751[79:64]     = Conv_out[65];
    assign  image_1_751[63:48]     = Conv_out[64];
    assign  image_1_751[47:32]     = Conv_out[36];
    assign  image_1_751[31:16]     = Conv_out[35];
    assign  image_1_751[15:0]      = Conv_out[34];

    assign  image_1_752[143:128]   = Conv_out[95];
    assign  image_1_752[127:112]   = Conv_out[94];
    assign  image_1_752[111:96]    = Conv_out[93];
    assign  image_1_752[95:80]     = Conv_out[65];
    assign  image_1_752[79:64]     = Conv_out[64];
    assign  image_1_752[63:48]     = Conv_out[63];
    assign  image_1_752[47:32]     = Conv_out[35];
    assign  image_1_752[31:16]     = Conv_out[34];
    assign  image_1_752[15:0]      = Conv_out[33];

    assign  image_1_753[143:128]   = Conv_out[94];
    assign  image_1_753[127:112]   = Conv_out[93];
    assign  image_1_753[111:96]    = Conv_out[92];
    assign  image_1_753[95:80]     = Conv_out[64];
    assign  image_1_753[79:64]     = Conv_out[63];
    assign  image_1_753[63:48]     = Conv_out[62];
    assign  image_1_753[47:32]     = Conv_out[34];
    assign  image_1_753[31:16]     = Conv_out[33];
    assign  image_1_753[15:0]      = Conv_out[32];

    assign  image_1_754[143:128]   = Conv_out[93];
    assign  image_1_754[127:112]   = Conv_out[92];
    assign  image_1_754[111:96]    = Conv_out[91];
    assign  image_1_754[95:80]     = Conv_out[63];
    assign  image_1_754[79:64]     = Conv_out[62];
    assign  image_1_754[63:48]     = Conv_out[61];
    assign  image_1_754[47:32]     = Conv_out[33];
    assign  image_1_754[31:16]     = Conv_out[32];
    assign  image_1_754[15:0]      = Conv_out[31];

    assign  image_1_755[143:128]   = Conv_out[92];
    assign  image_1_755[127:112]   = Conv_out[91];
    assign  image_1_755[111:96]    = Conv_out[90];
    assign  image_1_755[95:80]     = Conv_out[62];
    assign  image_1_755[79:64]     = Conv_out[61];
    assign  image_1_755[63:48]     = Conv_out[60];
    assign  image_1_755[47:32]     = Conv_out[32];
    assign  image_1_755[31:16]     = Conv_out[31];
    assign  image_1_755[15:0]      = Conv_out[30];

    assign  image_1_756[143:128]   = Conv_out[89];
    assign  image_1_756[127:112]   = Conv_out[88];
    assign  image_1_756[111:96]    = Conv_out[87];
    assign  image_1_756[95:80]     = Conv_out[59];
    assign  image_1_756[79:64]     = Conv_out[58];
    assign  image_1_756[63:48]     = Conv_out[57];
    assign  image_1_756[47:32]     = Conv_out[29];
    assign  image_1_756[31:16]     = Conv_out[28];
    assign  image_1_756[15:0]      = Conv_out[27];

    assign  image_1_757[143:128]   = Conv_out[88];
    assign  image_1_757[127:112]   = Conv_out[87];
    assign  image_1_757[111:96]    = Conv_out[86];
    assign  image_1_757[95:80]     = Conv_out[58];
    assign  image_1_757[79:64]     = Conv_out[57];
    assign  image_1_757[63:48]     = Conv_out[56];
    assign  image_1_757[47:32]     = Conv_out[28];
    assign  image_1_757[31:16]     = Conv_out[27];
    assign  image_1_757[15:0]      = Conv_out[26];

    assign  image_1_758[143:128]   = Conv_out[87];
    assign  image_1_758[127:112]   = Conv_out[86];
    assign  image_1_758[111:96]    = Conv_out[85];
    assign  image_1_758[95:80]     = Conv_out[57];
    assign  image_1_758[79:64]     = Conv_out[56];
    assign  image_1_758[63:48]     = Conv_out[55];
    assign  image_1_758[47:32]     = Conv_out[27];
    assign  image_1_758[31:16]     = Conv_out[26];
    assign  image_1_758[15:0]      = Conv_out[25];

    assign  image_1_759[143:128]   = Conv_out[86];
    assign  image_1_759[127:112]   = Conv_out[85];
    assign  image_1_759[111:96]    = Conv_out[84];
    assign  image_1_759[95:80]     = Conv_out[56];
    assign  image_1_759[79:64]     = Conv_out[55];
    assign  image_1_759[63:48]     = Conv_out[54];
    assign  image_1_759[47:32]     = Conv_out[26];
    assign  image_1_759[31:16]     = Conv_out[25];
    assign  image_1_759[15:0]      = Conv_out[24];

    assign  image_1_760[143:128]   = Conv_out[85];
    assign  image_1_760[127:112]   = Conv_out[84];
    assign  image_1_760[111:96]    = Conv_out[83];
    assign  image_1_760[95:80]     = Conv_out[55];
    assign  image_1_760[79:64]     = Conv_out[54];
    assign  image_1_760[63:48]     = Conv_out[53];
    assign  image_1_760[47:32]     = Conv_out[25];
    assign  image_1_760[31:16]     = Conv_out[24];
    assign  image_1_760[15:0]      = Conv_out[23];

    assign  image_1_761[143:128]   = Conv_out[84];
    assign  image_1_761[127:112]   = Conv_out[83];
    assign  image_1_761[111:96]    = Conv_out[82];
    assign  image_1_761[95:80]     = Conv_out[54];
    assign  image_1_761[79:64]     = Conv_out[53];
    assign  image_1_761[63:48]     = Conv_out[52];
    assign  image_1_761[47:32]     = Conv_out[24];
    assign  image_1_761[31:16]     = Conv_out[23];
    assign  image_1_761[15:0]      = Conv_out[22];

    assign  image_1_762[143:128]   = Conv_out[83];
    assign  image_1_762[127:112]   = Conv_out[82];
    assign  image_1_762[111:96]    = Conv_out[81];
    assign  image_1_762[95:80]     = Conv_out[53];
    assign  image_1_762[79:64]     = Conv_out[52];
    assign  image_1_762[63:48]     = Conv_out[51];
    assign  image_1_762[47:32]     = Conv_out[23];
    assign  image_1_762[31:16]     = Conv_out[22];
    assign  image_1_762[15:0]      = Conv_out[21];

    assign  image_1_763[143:128]   = Conv_out[82];
    assign  image_1_763[127:112]   = Conv_out[81];
    assign  image_1_763[111:96]    = Conv_out[80];
    assign  image_1_763[95:80]     = Conv_out[52];
    assign  image_1_763[79:64]     = Conv_out[51];
    assign  image_1_763[63:48]     = Conv_out[50];
    assign  image_1_763[47:32]     = Conv_out[22];
    assign  image_1_763[31:16]     = Conv_out[21];
    assign  image_1_763[15:0]      = Conv_out[20];

    assign  image_1_764[143:128]   = Conv_out[81];
    assign  image_1_764[127:112]   = Conv_out[80];
    assign  image_1_764[111:96]    = Conv_out[79];
    assign  image_1_764[95:80]     = Conv_out[51];
    assign  image_1_764[79:64]     = Conv_out[50];
    assign  image_1_764[63:48]     = Conv_out[49];
    assign  image_1_764[47:32]     = Conv_out[21];
    assign  image_1_764[31:16]     = Conv_out[20];
    assign  image_1_764[15:0]      = Conv_out[19];

    assign  image_1_765[143:128]   = Conv_out[80];
    assign  image_1_765[127:112]   = Conv_out[79];
    assign  image_1_765[111:96]    = Conv_out[78];
    assign  image_1_765[95:80]     = Conv_out[50];
    assign  image_1_765[79:64]     = Conv_out[49];
    assign  image_1_765[63:48]     = Conv_out[48];
    assign  image_1_765[47:32]     = Conv_out[20];
    assign  image_1_765[31:16]     = Conv_out[19];
    assign  image_1_765[15:0]      = Conv_out[18];

    assign  image_1_766[143:128]   = Conv_out[79];
    assign  image_1_766[127:112]   = Conv_out[78];
    assign  image_1_766[111:96]    = Conv_out[77];
    assign  image_1_766[95:80]     = Conv_out[49];
    assign  image_1_766[79:64]     = Conv_out[48];
    assign  image_1_766[63:48]     = Conv_out[47];
    assign  image_1_766[47:32]     = Conv_out[19];
    assign  image_1_766[31:16]     = Conv_out[18];
    assign  image_1_766[15:0]      = Conv_out[17];

    assign  image_1_767[143:128]   = Conv_out[78];
    assign  image_1_767[127:112]   = Conv_out[77];
    assign  image_1_767[111:96]    = Conv_out[76];
    assign  image_1_767[95:80]     = Conv_out[48];
    assign  image_1_767[79:64]     = Conv_out[47];
    assign  image_1_767[63:48]     = Conv_out[46];
    assign  image_1_767[47:32]     = Conv_out[18];
    assign  image_1_767[31:16]     = Conv_out[17];
    assign  image_1_767[15:0]      = Conv_out[16];

    assign  image_1_768[143:128]   = Conv_out[77];
    assign  image_1_768[127:112]   = Conv_out[76];
    assign  image_1_768[111:96]    = Conv_out[75];
    assign  image_1_768[95:80]     = Conv_out[47];
    assign  image_1_768[79:64]     = Conv_out[46];
    assign  image_1_768[63:48]     = Conv_out[45];
    assign  image_1_768[47:32]     = Conv_out[17];
    assign  image_1_768[31:16]     = Conv_out[16];
    assign  image_1_768[15:0]      = Conv_out[15];

    assign  image_1_769[143:128]   = Conv_out[76];
    assign  image_1_769[127:112]   = Conv_out[75];
    assign  image_1_769[111:96]    = Conv_out[74];
    assign  image_1_769[95:80]     = Conv_out[46];
    assign  image_1_769[79:64]     = Conv_out[45];
    assign  image_1_769[63:48]     = Conv_out[44];
    assign  image_1_769[47:32]     = Conv_out[16];
    assign  image_1_769[31:16]     = Conv_out[15];
    assign  image_1_769[15:0]      = Conv_out[14];

    assign  image_1_770[143:128]   = Conv_out[75];
    assign  image_1_770[127:112]   = Conv_out[74];
    assign  image_1_770[111:96]    = Conv_out[73];
    assign  image_1_770[95:80]     = Conv_out[45];
    assign  image_1_770[79:64]     = Conv_out[44];
    assign  image_1_770[63:48]     = Conv_out[43];
    assign  image_1_770[47:32]     = Conv_out[15];
    assign  image_1_770[31:16]     = Conv_out[14];
    assign  image_1_770[15:0]      = Conv_out[13];

    assign  image_1_771[143:128]   = Conv_out[74];
    assign  image_1_771[127:112]   = Conv_out[73];
    assign  image_1_771[111:96]    = Conv_out[72];
    assign  image_1_771[95:80]     = Conv_out[44];
    assign  image_1_771[79:64]     = Conv_out[43];
    assign  image_1_771[63:48]     = Conv_out[42];
    assign  image_1_771[47:32]     = Conv_out[14];
    assign  image_1_771[31:16]     = Conv_out[13];
    assign  image_1_771[15:0]      = Conv_out[12];

    assign  image_1_772[143:128]   = Conv_out[73];
    assign  image_1_772[127:112]   = Conv_out[72];
    assign  image_1_772[111:96]    = Conv_out[71];
    assign  image_1_772[95:80]     = Conv_out[43];
    assign  image_1_772[79:64]     = Conv_out[42];
    assign  image_1_772[63:48]     = Conv_out[41];
    assign  image_1_772[47:32]     = Conv_out[13];
    assign  image_1_772[31:16]     = Conv_out[12];
    assign  image_1_772[15:0]      = Conv_out[11];

    assign  image_1_773[143:128]   = Conv_out[72];
    assign  image_1_773[127:112]   = Conv_out[71];
    assign  image_1_773[111:96]    = Conv_out[70];
    assign  image_1_773[95:80]     = Conv_out[42];
    assign  image_1_773[79:64]     = Conv_out[41];
    assign  image_1_773[63:48]     = Conv_out[40];
    assign  image_1_773[47:32]     = Conv_out[12];
    assign  image_1_773[31:16]     = Conv_out[11];
    assign  image_1_773[15:0]      = Conv_out[10];

    assign  image_1_774[143:128]   = Conv_out[71];
    assign  image_1_774[127:112]   = Conv_out[70];
    assign  image_1_774[111:96]    = Conv_out[69];
    assign  image_1_774[95:80]     = Conv_out[41];
    assign  image_1_774[79:64]     = Conv_out[40];
    assign  image_1_774[63:48]     = Conv_out[39];
    assign  image_1_774[47:32]     = Conv_out[11];
    assign  image_1_774[31:16]     = Conv_out[10];
    assign  image_1_774[15:0]      = Conv_out[9];

    assign  image_1_775[143:128]   = Conv_out[70];
    assign  image_1_775[127:112]   = Conv_out[69];
    assign  image_1_775[111:96]    = Conv_out[68];
    assign  image_1_775[95:80]     = Conv_out[40];
    assign  image_1_775[79:64]     = Conv_out[39];
    assign  image_1_775[63:48]     = Conv_out[38];
    assign  image_1_775[47:32]     = Conv_out[10];
    assign  image_1_775[31:16]     = Conv_out[9];
    assign  image_1_775[15:0]      = Conv_out[8];

    assign  image_1_776[143:128]   = Conv_out[69];
    assign  image_1_776[127:112]   = Conv_out[68];
    assign  image_1_776[111:96]    = Conv_out[67];
    assign  image_1_776[95:80]     = Conv_out[39];
    assign  image_1_776[79:64]     = Conv_out[38];
    assign  image_1_776[63:48]     = Conv_out[37];
    assign  image_1_776[47:32]     = Conv_out[9];
    assign  image_1_776[31:16]     = Conv_out[8];
    assign  image_1_776[15:0]      = Conv_out[7];

    assign  image_1_777[143:128]   = Conv_out[68];
    assign  image_1_777[127:112]   = Conv_out[67];
    assign  image_1_777[111:96]    = Conv_out[66];
    assign  image_1_777[95:80]     = Conv_out[38];
    assign  image_1_777[79:64]     = Conv_out[37];
    assign  image_1_777[63:48]     = Conv_out[36];
    assign  image_1_777[47:32]     = Conv_out[8];
    assign  image_1_777[31:16]     = Conv_out[7];
    assign  image_1_777[15:0]      = Conv_out[6];

    assign  image_1_778[143:128]   = Conv_out[67];
    assign  image_1_778[127:112]   = Conv_out[66];
    assign  image_1_778[111:96]    = Conv_out[65];
    assign  image_1_778[95:80]     = Conv_out[37];
    assign  image_1_778[79:64]     = Conv_out[36];
    assign  image_1_778[63:48]     = Conv_out[35];
    assign  image_1_778[47:32]     = Conv_out[7];
    assign  image_1_778[31:16]     = Conv_out[6];
    assign  image_1_778[15:0]      = Conv_out[5];

    assign  image_1_779[143:128]   = Conv_out[66];
    assign  image_1_779[127:112]   = Conv_out[65];
    assign  image_1_779[111:96]    = Conv_out[64];
    assign  image_1_779[95:80]     = Conv_out[36];
    assign  image_1_779[79:64]     = Conv_out[35];
    assign  image_1_779[63:48]     = Conv_out[34];
    assign  image_1_779[47:32]     = Conv_out[6];
    assign  image_1_779[31:16]     = Conv_out[5];
    assign  image_1_779[15:0]      = Conv_out[4];

    assign  image_1_780[143:128]   = Conv_out[65];
    assign  image_1_780[127:112]   = Conv_out[64];
    assign  image_1_780[111:96]    = Conv_out[63];
    assign  image_1_780[95:80]     = Conv_out[35];
    assign  image_1_780[79:64]     = Conv_out[34];
    assign  image_1_780[63:48]     = Conv_out[33];
    assign  image_1_780[47:32]     = Conv_out[5];
    assign  image_1_780[31:16]     = Conv_out[4];
    assign  image_1_780[15:0]      = Conv_out[3];

    assign  image_1_781[143:128]   = Conv_out[64];
    assign  image_1_781[127:112]   = Conv_out[63];
    assign  image_1_781[111:96]    = Conv_out[62];
    assign  image_1_781[95:80]     = Conv_out[34];
    assign  image_1_781[79:64]     = Conv_out[33];
    assign  image_1_781[63:48]     = Conv_out[32];
    assign  image_1_781[47:32]     = Conv_out[4];
    assign  image_1_781[31:16]     = Conv_out[3];
    assign  image_1_781[15:0]      = Conv_out[2];

    assign  image_1_782[143:128]   = Conv_out[63];
    assign  image_1_782[127:112]   = Conv_out[62];
    assign  image_1_782[111:96]    = Conv_out[61];
    assign  image_1_782[95:80]     = Conv_out[33];
    assign  image_1_782[79:64]     = Conv_out[32];
    assign  image_1_782[63:48]     = Conv_out[31];
    assign  image_1_782[47:32]     = Conv_out[3];
    assign  image_1_782[31:16]     = Conv_out[2];
    assign  image_1_782[15:0]      = Conv_out[1];

    assign  image_1_783[143:128]   = Conv_out[62];
    assign  image_1_783[127:112]   = Conv_out[61];
    assign  image_1_783[111:96]    = Conv_out[60];
    assign  image_1_783[95:80]     = Conv_out[32];
    assign  image_1_783[79:64]     = Conv_out[31];
    assign  image_1_783[63:48]     = Conv_out[30];
    assign  image_1_783[47:32]     = Conv_out[2];
    assign  image_1_783[31:16]     = Conv_out[1];
    assign  image_1_783[15:0]      = Conv_out[0];


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
CNN_Single_Layer    single_0(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_0), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_899)
    );

CNN_Single_Layer    single_1(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_1), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_898)
    );

CNN_Single_Layer    single_2(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_2), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_897)
    );

CNN_Single_Layer    single_3(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_3), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_896)
    );

CNN_Single_Layer    single_4(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_4), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_895)
    );

CNN_Single_Layer    single_5(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_5), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_894)
    );

CNN_Single_Layer    single_6(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_6), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_893)
    );

CNN_Single_Layer    single_7(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_7), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_892)
    );

CNN_Single_Layer    single_8(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_8), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_891)
    );

CNN_Single_Layer    single_9(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_9), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_890)
    );

CNN_Single_Layer    single_10(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_10), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_889)
    );

CNN_Single_Layer    single_11(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_11), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_888)
    );

CNN_Single_Layer    single_12(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_12), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_887)
    );

CNN_Single_Layer    single_13(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_13), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_886)
    );

CNN_Single_Layer    single_14(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_14), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_885)
    );

CNN_Single_Layer    single_15(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_15), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_884)
    );

CNN_Single_Layer    single_16(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_16), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_883)
    );

CNN_Single_Layer    single_17(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_17), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_882)
    );

CNN_Single_Layer    single_18(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_18), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_881)
    );

CNN_Single_Layer    single_19(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_19), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_880)
    );

CNN_Single_Layer    single_20(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_20), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_879)
    );

CNN_Single_Layer    single_21(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_21), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_878)
    );

CNN_Single_Layer    single_22(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_22), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_877)
    );

CNN_Single_Layer    single_23(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_23), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_876)
    );

CNN_Single_Layer    single_24(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_24), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_875)
    );

CNN_Single_Layer    single_25(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_25), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_874)
    );

CNN_Single_Layer    single_26(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_26), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_873)
    );

CNN_Single_Layer    single_27(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_27), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_872)
    );

CNN_Single_Layer    single_28(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_28), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_871)
    );

CNN_Single_Layer    single_29(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_29), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_870)
    );

CNN_Single_Layer    single_30(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_30), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_869)
    );

CNN_Single_Layer    single_31(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_31), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_868)
    );

CNN_Single_Layer    single_32(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_32), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_867)
    );

CNN_Single_Layer    single_33(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_33), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_866)
    );

CNN_Single_Layer    single_34(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_34), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_865)
    );

CNN_Single_Layer    single_35(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_35), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_864)
    );

CNN_Single_Layer    single_36(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_36), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_863)
    );

CNN_Single_Layer    single_37(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_37), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_862)
    );

CNN_Single_Layer    single_38(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_38), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_861)
    );

CNN_Single_Layer    single_39(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_39), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_860)
    );

CNN_Single_Layer    single_40(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_40), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_859)
    );

CNN_Single_Layer    single_41(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_41), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_858)
    );

CNN_Single_Layer    single_42(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_42), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_857)
    );

CNN_Single_Layer    single_43(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_43), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_856)
    );

CNN_Single_Layer    single_44(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_44), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_855)
    );

CNN_Single_Layer    single_45(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_45), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_854)
    );

CNN_Single_Layer    single_46(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_46), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_853)
    );

CNN_Single_Layer    single_47(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_47), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_852)
    );

CNN_Single_Layer    single_48(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_48), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_851)
    );

CNN_Single_Layer    single_49(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_49), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_850)
    );

CNN_Single_Layer    single_50(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_50), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_849)
    );

CNN_Single_Layer    single_51(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_51), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_848)
    );

CNN_Single_Layer    single_52(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_52), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_847)
    );

CNN_Single_Layer    single_53(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_53), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_846)
    );

CNN_Single_Layer    single_54(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_54), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_845)
    );

CNN_Single_Layer    single_55(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_55), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_844)
    );

CNN_Single_Layer    single_56(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_56), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_843)
    );

CNN_Single_Layer    single_57(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_57), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_842)
    );

CNN_Single_Layer    single_58(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_58), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_841)
    );

CNN_Single_Layer    single_59(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_59), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_840)
    );

CNN_Single_Layer    single_60(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_60), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_839)
    );

CNN_Single_Layer    single_61(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_61), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_838)
    );

CNN_Single_Layer    single_62(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_62), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_837)
    );

CNN_Single_Layer    single_63(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_63), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_836)
    );

CNN_Single_Layer    single_64(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_64), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_835)
    );

CNN_Single_Layer    single_65(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_65), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_834)
    );

CNN_Single_Layer    single_66(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_66), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_833)
    );

CNN_Single_Layer    single_67(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_67), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_832)
    );

CNN_Single_Layer    single_68(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_68), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_831)
    );

CNN_Single_Layer    single_69(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_69), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_830)
    );

CNN_Single_Layer    single_70(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_70), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_829)
    );

CNN_Single_Layer    single_71(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_71), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_828)
    );

CNN_Single_Layer    single_72(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_72), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_827)
    );

CNN_Single_Layer    single_73(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_73), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_826)
    );

CNN_Single_Layer    single_74(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_74), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_825)
    );

CNN_Single_Layer    single_75(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_75), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_824)
    );

CNN_Single_Layer    single_76(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_76), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_823)
    );

CNN_Single_Layer    single_77(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_77), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_822)
    );

CNN_Single_Layer    single_78(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_78), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_821)
    );

CNN_Single_Layer    single_79(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_79), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_820)
    );

CNN_Single_Layer    single_80(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_80), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_819)
    );

CNN_Single_Layer    single_81(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_81), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_818)
    );

CNN_Single_Layer    single_82(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_82), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_817)
    );

CNN_Single_Layer    single_83(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_83), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_816)
    );

CNN_Single_Layer    single_84(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_84), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_815)
    );

CNN_Single_Layer    single_85(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_85), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_814)
    );

CNN_Single_Layer    single_86(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_86), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_813)
    );

CNN_Single_Layer    single_87(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_87), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_812)
    );

CNN_Single_Layer    single_88(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_88), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_811)
    );

CNN_Single_Layer    single_89(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_89), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_810)
    );

CNN_Single_Layer    single_90(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_90), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_809)
    );

CNN_Single_Layer    single_91(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_91), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_808)
    );

CNN_Single_Layer    single_92(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_92), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_807)
    );

CNN_Single_Layer    single_93(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_93), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_806)
    );

CNN_Single_Layer    single_94(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_94), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_805)
    );

CNN_Single_Layer    single_95(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_95), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_804)
    );

CNN_Single_Layer    single_96(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_96), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_803)
    );

CNN_Single_Layer    single_97(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_97), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_802)
    );

CNN_Single_Layer    single_98(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_98), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_801)
    );

CNN_Single_Layer    single_99(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_99), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_800)
    );

CNN_Single_Layer    single_100(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_100), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_799)
    );

CNN_Single_Layer    single_101(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_101), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_798)
    );

CNN_Single_Layer    single_102(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_102), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_797)
    );

CNN_Single_Layer    single_103(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_103), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_796)
    );

CNN_Single_Layer    single_104(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_104), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_795)
    );

CNN_Single_Layer    single_105(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_105), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_794)
    );

CNN_Single_Layer    single_106(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_106), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_793)
    );

CNN_Single_Layer    single_107(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_107), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_792)
    );

CNN_Single_Layer    single_108(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_108), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_791)
    );

CNN_Single_Layer    single_109(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_109), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_790)
    );

CNN_Single_Layer    single_110(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_110), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_789)
    );

CNN_Single_Layer    single_111(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_111), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_788)
    );

CNN_Single_Layer    single_112(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_112), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_787)
    );

CNN_Single_Layer    single_113(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_113), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_786)
    );

CNN_Single_Layer    single_114(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_114), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_785)
    );

CNN_Single_Layer    single_115(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_115), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_784)
    );

CNN_Single_Layer    single_116(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_116), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_783)
    );

CNN_Single_Layer    single_117(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_117), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_782)
    );

CNN_Single_Layer    single_118(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_118), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_781)
    );

CNN_Single_Layer    single_119(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_119), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_780)
    );

CNN_Single_Layer    single_120(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_120), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_779)
    );

CNN_Single_Layer    single_121(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_121), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_778)
    );

CNN_Single_Layer    single_122(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_122), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_777)
    );

CNN_Single_Layer    single_123(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_123), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_776)
    );

CNN_Single_Layer    single_124(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_124), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_775)
    );

CNN_Single_Layer    single_125(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_125), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_774)
    );

CNN_Single_Layer    single_126(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_126), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_773)
    );

CNN_Single_Layer    single_127(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_127), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_772)
    );

CNN_Single_Layer    single_128(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_128), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_771)
    );

CNN_Single_Layer    single_129(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_129), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_770)
    );

CNN_Single_Layer    single_130(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_130), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_769)
    );

CNN_Single_Layer    single_131(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_131), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_768)
    );

CNN_Single_Layer    single_132(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_132), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_767)
    );

CNN_Single_Layer    single_133(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_133), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_766)
    );

CNN_Single_Layer    single_134(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_134), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_765)
    );

CNN_Single_Layer    single_135(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_135), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_764)
    );

CNN_Single_Layer    single_136(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_136), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_763)
    );

CNN_Single_Layer    single_137(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_137), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_762)
    );

CNN_Single_Layer    single_138(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_138), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_761)
    );

CNN_Single_Layer    single_139(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_139), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_760)
    );

CNN_Single_Layer    single_140(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_140), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_759)
    );

CNN_Single_Layer    single_141(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_141), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_758)
    );

CNN_Single_Layer    single_142(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_142), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_757)
    );

CNN_Single_Layer    single_143(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_143), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_756)
    );

CNN_Single_Layer    single_144(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_144), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_755)
    );

CNN_Single_Layer    single_145(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_145), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_754)
    );

CNN_Single_Layer    single_146(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_146), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_753)
    );

CNN_Single_Layer    single_147(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_147), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_752)
    );

CNN_Single_Layer    single_148(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_148), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_751)
    );

CNN_Single_Layer    single_149(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_149), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_750)
    );

CNN_Single_Layer    single_150(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_150), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_749)
    );

CNN_Single_Layer    single_151(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_151), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_748)
    );

CNN_Single_Layer    single_152(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_152), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_747)
    );

CNN_Single_Layer    single_153(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_153), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_746)
    );

CNN_Single_Layer    single_154(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_154), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_745)
    );

CNN_Single_Layer    single_155(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_155), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_744)
    );

CNN_Single_Layer    single_156(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_156), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_743)
    );

CNN_Single_Layer    single_157(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_157), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_742)
    );

CNN_Single_Layer    single_158(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_158), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_741)
    );

CNN_Single_Layer    single_159(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_159), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_740)
    );

CNN_Single_Layer    single_160(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_160), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_739)
    );

CNN_Single_Layer    single_161(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_161), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_738)
    );

CNN_Single_Layer    single_162(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_162), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_737)
    );

CNN_Single_Layer    single_163(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_163), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_736)
    );

CNN_Single_Layer    single_164(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_164), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_735)
    );

CNN_Single_Layer    single_165(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_165), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_734)
    );

CNN_Single_Layer    single_166(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_166), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_733)
    );

CNN_Single_Layer    single_167(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_167), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_732)
    );

CNN_Single_Layer    single_168(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_168), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_731)
    );

CNN_Single_Layer    single_169(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_169), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_730)
    );

CNN_Single_Layer    single_170(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_170), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_729)
    );

CNN_Single_Layer    single_171(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_171), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_728)
    );

CNN_Single_Layer    single_172(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_172), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_727)
    );

CNN_Single_Layer    single_173(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_173), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_726)
    );

CNN_Single_Layer    single_174(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_174), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_725)
    );

CNN_Single_Layer    single_175(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_175), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_724)
    );

CNN_Single_Layer    single_176(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_176), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_723)
    );

CNN_Single_Layer    single_177(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_177), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_722)
    );

CNN_Single_Layer    single_178(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_178), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_721)
    );

CNN_Single_Layer    single_179(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_179), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_720)
    );

CNN_Single_Layer    single_180(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_180), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_719)
    );

CNN_Single_Layer    single_181(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_181), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_718)
    );

CNN_Single_Layer    single_182(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_182), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_717)
    );

CNN_Single_Layer    single_183(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_183), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_716)
    );

CNN_Single_Layer    single_184(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_184), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_715)
    );

CNN_Single_Layer    single_185(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_185), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_714)
    );

CNN_Single_Layer    single_186(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_186), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_713)
    );

CNN_Single_Layer    single_187(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_187), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_712)
    );

CNN_Single_Layer    single_188(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_188), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_711)
    );

CNN_Single_Layer    single_189(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_189), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_710)
    );

CNN_Single_Layer    single_190(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_190), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_709)
    );

CNN_Single_Layer    single_191(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_191), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_708)
    );

CNN_Single_Layer    single_192(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_192), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_707)
    );

CNN_Single_Layer    single_193(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_193), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_706)
    );

CNN_Single_Layer    single_194(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_194), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_705)
    );

CNN_Single_Layer    single_195(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_195), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_704)
    );

CNN_Single_Layer    single_196(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_196), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_703)
    );

CNN_Single_Layer    single_197(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_197), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_702)
    );

CNN_Single_Layer    single_198(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_198), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_701)
    );

CNN_Single_Layer    single_199(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_199), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_700)
    );

CNN_Single_Layer    single_200(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_200), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_699)
    );

CNN_Single_Layer    single_201(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_201), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_698)
    );

CNN_Single_Layer    single_202(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_202), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_697)
    );

CNN_Single_Layer    single_203(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_203), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_696)
    );

CNN_Single_Layer    single_204(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_204), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_695)
    );

CNN_Single_Layer    single_205(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_205), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_694)
    );

CNN_Single_Layer    single_206(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_206), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_693)
    );

CNN_Single_Layer    single_207(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_207), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_692)
    );

CNN_Single_Layer    single_208(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_208), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_691)
    );

CNN_Single_Layer    single_209(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_209), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_690)
    );

CNN_Single_Layer    single_210(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_210), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_689)
    );

CNN_Single_Layer    single_211(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_211), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_688)
    );

CNN_Single_Layer    single_212(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_212), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_687)
    );

CNN_Single_Layer    single_213(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_213), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_686)
    );

CNN_Single_Layer    single_214(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_214), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_685)
    );

CNN_Single_Layer    single_215(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_215), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_684)
    );

CNN_Single_Layer    single_216(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_216), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_683)
    );

CNN_Single_Layer    single_217(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_217), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_682)
    );

CNN_Single_Layer    single_218(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_218), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_681)
    );

CNN_Single_Layer    single_219(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_219), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_680)
    );

CNN_Single_Layer    single_220(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_220), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_679)
    );

CNN_Single_Layer    single_221(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_221), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_678)
    );

CNN_Single_Layer    single_222(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_222), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_677)
    );

CNN_Single_Layer    single_223(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_223), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_676)
    );

CNN_Single_Layer    single_224(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_224), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_675)
    );

CNN_Single_Layer    single_225(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_225), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_674)
    );

CNN_Single_Layer    single_226(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_226), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_673)
    );

CNN_Single_Layer    single_227(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_227), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_672)
    );

CNN_Single_Layer    single_228(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_228), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_671)
    );

CNN_Single_Layer    single_229(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_229), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_670)
    );

CNN_Single_Layer    single_230(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_230), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_669)
    );

CNN_Single_Layer    single_231(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_231), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_668)
    );

CNN_Single_Layer    single_232(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_232), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_667)
    );

CNN_Single_Layer    single_233(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_233), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_666)
    );

CNN_Single_Layer    single_234(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_234), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_665)
    );

CNN_Single_Layer    single_235(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_235), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_664)
    );

CNN_Single_Layer    single_236(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_236), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_663)
    );

CNN_Single_Layer    single_237(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_237), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_662)
    );

CNN_Single_Layer    single_238(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_238), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_661)
    );

CNN_Single_Layer    single_239(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_239), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_660)
    );

CNN_Single_Layer    single_240(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_240), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_659)
    );

CNN_Single_Layer    single_241(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_241), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_658)
    );

CNN_Single_Layer    single_242(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_242), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_657)
    );

CNN_Single_Layer    single_243(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_243), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_656)
    );

CNN_Single_Layer    single_244(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_244), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_655)
    );

CNN_Single_Layer    single_245(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_245), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_654)
    );

CNN_Single_Layer    single_246(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_246), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_653)
    );

CNN_Single_Layer    single_247(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_247), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_652)
    );

CNN_Single_Layer    single_248(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_248), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_651)
    );

CNN_Single_Layer    single_249(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_249), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_650)
    );

CNN_Single_Layer    single_250(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_250), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_649)
    );

CNN_Single_Layer    single_251(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_251), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_648)
    );

CNN_Single_Layer    single_252(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_252), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_647)
    );

CNN_Single_Layer    single_253(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_253), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_646)
    );

CNN_Single_Layer    single_254(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_254), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_645)
    );

CNN_Single_Layer    single_255(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_255), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_644)
    );

CNN_Single_Layer    single_256(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_256), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_643)
    );

CNN_Single_Layer    single_257(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_257), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_642)
    );

CNN_Single_Layer    single_258(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_258), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_641)
    );

CNN_Single_Layer    single_259(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_259), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_640)
    );

CNN_Single_Layer    single_260(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_260), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_639)
    );

CNN_Single_Layer    single_261(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_261), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_638)
    );

CNN_Single_Layer    single_262(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_262), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_637)
    );

CNN_Single_Layer    single_263(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_263), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_636)
    );

CNN_Single_Layer    single_264(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_264), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_635)
    );

CNN_Single_Layer    single_265(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_265), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_634)
    );

CNN_Single_Layer    single_266(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_266), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_633)
    );

CNN_Single_Layer    single_267(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_267), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_632)
    );

CNN_Single_Layer    single_268(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_268), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_631)
    );

CNN_Single_Layer    single_269(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_269), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_630)
    );

CNN_Single_Layer    single_270(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_270), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_629)
    );

CNN_Single_Layer    single_271(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_271), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_628)
    );

CNN_Single_Layer    single_272(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_272), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_627)
    );

CNN_Single_Layer    single_273(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_273), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_626)
    );

CNN_Single_Layer    single_274(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_274), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_625)
    );

CNN_Single_Layer    single_275(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_275), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_624)
    );

CNN_Single_Layer    single_276(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_276), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_623)
    );

CNN_Single_Layer    single_277(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_277), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_622)
    );

CNN_Single_Layer    single_278(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_278), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_621)
    );

CNN_Single_Layer    single_279(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_279), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_620)
    );

CNN_Single_Layer    single_280(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_280), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_619)
    );

CNN_Single_Layer    single_281(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_281), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_618)
    );

CNN_Single_Layer    single_282(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_282), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_617)
    );

CNN_Single_Layer    single_283(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_283), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_616)
    );

CNN_Single_Layer    single_284(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_284), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_615)
    );

CNN_Single_Layer    single_285(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_285), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_614)
    );

CNN_Single_Layer    single_286(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_286), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_613)
    );

CNN_Single_Layer    single_287(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_287), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_612)
    );

CNN_Single_Layer    single_288(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_288), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_611)
    );

CNN_Single_Layer    single_289(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_289), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_610)
    );

CNN_Single_Layer    single_290(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_290), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_609)
    );

CNN_Single_Layer    single_291(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_291), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_608)
    );

CNN_Single_Layer    single_292(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_292), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_607)
    );

CNN_Single_Layer    single_293(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_293), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_606)
    );

CNN_Single_Layer    single_294(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_294), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_605)
    );

CNN_Single_Layer    single_295(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_295), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_604)
    );

CNN_Single_Layer    single_296(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_296), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_603)
    );

CNN_Single_Layer    single_297(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_297), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_602)
    );

CNN_Single_Layer    single_298(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_298), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_601)
    );

CNN_Single_Layer    single_299(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_299), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_600)
    );

CNN_Single_Layer    single_300(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_300), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_599)
    );

CNN_Single_Layer    single_301(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_301), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_598)
    );

CNN_Single_Layer    single_302(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_302), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_597)
    );

CNN_Single_Layer    single_303(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_303), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_596)
    );

CNN_Single_Layer    single_304(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_304), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_595)
    );

CNN_Single_Layer    single_305(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_305), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_594)
    );

CNN_Single_Layer    single_306(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_306), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_593)
    );

CNN_Single_Layer    single_307(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_307), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_592)
    );

CNN_Single_Layer    single_308(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_308), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_591)
    );

CNN_Single_Layer    single_309(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_309), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_590)
    );

CNN_Single_Layer    single_310(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_310), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_589)
    );

CNN_Single_Layer    single_311(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_311), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_588)
    );

CNN_Single_Layer    single_312(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_312), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_587)
    );

CNN_Single_Layer    single_313(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_313), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_586)
    );

CNN_Single_Layer    single_314(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_314), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_585)
    );

CNN_Single_Layer    single_315(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_315), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_584)
    );

CNN_Single_Layer    single_316(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_316), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_583)
    );

CNN_Single_Layer    single_317(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_317), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_582)
    );

CNN_Single_Layer    single_318(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_318), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_581)
    );

CNN_Single_Layer    single_319(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_319), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_580)
    );

CNN_Single_Layer    single_320(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_320), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_579)
    );

CNN_Single_Layer    single_321(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_321), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_578)
    );

CNN_Single_Layer    single_322(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_322), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_577)
    );

CNN_Single_Layer    single_323(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_323), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_576)
    );

CNN_Single_Layer    single_324(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_324), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_575)
    );

CNN_Single_Layer    single_325(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_325), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_574)
    );

CNN_Single_Layer    single_326(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_326), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_573)
    );

CNN_Single_Layer    single_327(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_327), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_572)
    );

CNN_Single_Layer    single_328(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_328), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_571)
    );

CNN_Single_Layer    single_329(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_329), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_570)
    );

CNN_Single_Layer    single_330(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_330), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_569)
    );

CNN_Single_Layer    single_331(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_331), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_568)
    );

CNN_Single_Layer    single_332(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_332), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_567)
    );

CNN_Single_Layer    single_333(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_333), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_566)
    );

CNN_Single_Layer    single_334(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_334), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_565)
    );

CNN_Single_Layer    single_335(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_335), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_564)
    );

CNN_Single_Layer    single_336(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_336), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_563)
    );

CNN_Single_Layer    single_337(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_337), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_562)
    );

CNN_Single_Layer    single_338(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_338), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_561)
    );

CNN_Single_Layer    single_339(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_339), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_560)
    );

CNN_Single_Layer    single_340(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_340), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_559)
    );

CNN_Single_Layer    single_341(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_341), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_558)
    );

CNN_Single_Layer    single_342(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_342), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_557)
    );

CNN_Single_Layer    single_343(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_343), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_556)
    );

CNN_Single_Layer    single_344(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_344), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_555)
    );

CNN_Single_Layer    single_345(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_345), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_554)
    );

CNN_Single_Layer    single_346(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_346), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_553)
    );

CNN_Single_Layer    single_347(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_347), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_552)
    );

CNN_Single_Layer    single_348(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_348), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_551)
    );

CNN_Single_Layer    single_349(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_349), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_550)
    );

CNN_Single_Layer    single_350(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_350), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_549)
    );

CNN_Single_Layer    single_351(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_351), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_548)
    );

CNN_Single_Layer    single_352(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_352), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_547)
    );

CNN_Single_Layer    single_353(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_353), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_546)
    );

CNN_Single_Layer    single_354(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_354), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_545)
    );

CNN_Single_Layer    single_355(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_355), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_544)
    );

CNN_Single_Layer    single_356(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_356), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_543)
    );

CNN_Single_Layer    single_357(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_357), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_542)
    );

CNN_Single_Layer    single_358(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_358), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_541)
    );

CNN_Single_Layer    single_359(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_359), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_540)
    );

CNN_Single_Layer    single_360(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_360), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_539)
    );

CNN_Single_Layer    single_361(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_361), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_538)
    );

CNN_Single_Layer    single_362(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_362), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_537)
    );

CNN_Single_Layer    single_363(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_363), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_536)
    );

CNN_Single_Layer    single_364(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_364), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_535)
    );

CNN_Single_Layer    single_365(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_365), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_534)
    );

CNN_Single_Layer    single_366(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_366), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_533)
    );

CNN_Single_Layer    single_367(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_367), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_532)
    );

CNN_Single_Layer    single_368(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_368), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_531)
    );

CNN_Single_Layer    single_369(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_369), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_530)
    );

CNN_Single_Layer    single_370(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_370), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_529)
    );

CNN_Single_Layer    single_371(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_371), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_528)
    );

CNN_Single_Layer    single_372(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_372), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_527)
    );

CNN_Single_Layer    single_373(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_373), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_526)
    );

CNN_Single_Layer    single_374(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_374), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_525)
    );

CNN_Single_Layer    single_375(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_375), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_524)
    );

CNN_Single_Layer    single_376(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_376), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_523)
    );

CNN_Single_Layer    single_377(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_377), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_522)
    );

CNN_Single_Layer    single_378(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_378), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_521)
    );

CNN_Single_Layer    single_379(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_379), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_520)
    );

CNN_Single_Layer    single_380(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_380), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_519)
    );

CNN_Single_Layer    single_381(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_381), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_518)
    );

CNN_Single_Layer    single_382(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_382), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_517)
    );

CNN_Single_Layer    single_383(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_383), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_516)
    );

CNN_Single_Layer    single_384(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_384), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_515)
    );

CNN_Single_Layer    single_385(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_385), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_514)
    );

CNN_Single_Layer    single_386(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_386), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_513)
    );

CNN_Single_Layer    single_387(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_387), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_512)
    );

CNN_Single_Layer    single_388(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_388), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_511)
    );

CNN_Single_Layer    single_389(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_389), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_510)
    );

CNN_Single_Layer    single_390(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_390), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_509)
    );

CNN_Single_Layer    single_391(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_391), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_508)
    );

CNN_Single_Layer    single_392(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_392), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_507)
    );

CNN_Single_Layer    single_393(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_393), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_506)
    );

CNN_Single_Layer    single_394(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_394), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_505)
    );

CNN_Single_Layer    single_395(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_395), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_504)
    );

CNN_Single_Layer    single_396(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_396), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_503)
    );

CNN_Single_Layer    single_397(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_397), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_502)
    );

CNN_Single_Layer    single_398(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_398), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_501)
    );

CNN_Single_Layer    single_399(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_399), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_500)
    );

CNN_Single_Layer    single_400(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_400), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_499)
    );

CNN_Single_Layer    single_401(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_401), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_498)
    );

CNN_Single_Layer    single_402(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_402), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_497)
    );

CNN_Single_Layer    single_403(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_403), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_496)
    );

CNN_Single_Layer    single_404(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_404), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_495)
    );

CNN_Single_Layer    single_405(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_405), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_494)
    );

CNN_Single_Layer    single_406(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_406), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_493)
    );

CNN_Single_Layer    single_407(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_407), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_492)
    );

CNN_Single_Layer    single_408(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_408), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_491)
    );

CNN_Single_Layer    single_409(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_409), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_490)
    );

CNN_Single_Layer    single_410(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_410), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_489)
    );

CNN_Single_Layer    single_411(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_411), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_488)
    );

CNN_Single_Layer    single_412(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_412), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_487)
    );

CNN_Single_Layer    single_413(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_413), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_486)
    );

CNN_Single_Layer    single_414(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_414), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_485)
    );

CNN_Single_Layer    single_415(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_415), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_484)
    );

CNN_Single_Layer    single_416(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_416), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_483)
    );

CNN_Single_Layer    single_417(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_417), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_482)
    );

CNN_Single_Layer    single_418(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_418), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_481)
    );

CNN_Single_Layer    single_419(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_419), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_480)
    );

CNN_Single_Layer    single_420(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_420), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_479)
    );

CNN_Single_Layer    single_421(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_421), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_478)
    );

CNN_Single_Layer    single_422(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_422), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_477)
    );

CNN_Single_Layer    single_423(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_423), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_476)
    );

CNN_Single_Layer    single_424(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_424), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_475)
    );

CNN_Single_Layer    single_425(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_425), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_474)
    );

CNN_Single_Layer    single_426(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_426), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_473)
    );

CNN_Single_Layer    single_427(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_427), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_472)
    );

CNN_Single_Layer    single_428(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_428), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_471)
    );

CNN_Single_Layer    single_429(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_429), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_470)
    );

CNN_Single_Layer    single_430(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_430), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_469)
    );

CNN_Single_Layer    single_431(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_431), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_468)
    );

CNN_Single_Layer    single_432(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_432), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_467)
    );

CNN_Single_Layer    single_433(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_433), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_466)
    );

CNN_Single_Layer    single_434(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_434), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_465)
    );

CNN_Single_Layer    single_435(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_435), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_464)
    );

CNN_Single_Layer    single_436(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_436), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_463)
    );

CNN_Single_Layer    single_437(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_437), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_462)
    );

CNN_Single_Layer    single_438(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_438), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_461)
    );

CNN_Single_Layer    single_439(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_439), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_460)
    );

CNN_Single_Layer    single_440(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_440), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_459)
    );

CNN_Single_Layer    single_441(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_441), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_458)
    );

CNN_Single_Layer    single_442(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_442), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_457)
    );

CNN_Single_Layer    single_443(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_443), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_456)
    );

CNN_Single_Layer    single_444(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_444), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_455)
    );

CNN_Single_Layer    single_445(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_445), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_454)
    );

CNN_Single_Layer    single_446(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_446), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_453)
    );

CNN_Single_Layer    single_447(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_447), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_452)
    );

CNN_Single_Layer    single_448(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_448), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_451)
    );

CNN_Single_Layer    single_449(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_449), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_450)
    );

CNN_Single_Layer    single_450(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_450), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_449)
    );

CNN_Single_Layer    single_451(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_451), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_448)
    );

CNN_Single_Layer    single_452(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_452), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_447)
    );

CNN_Single_Layer    single_453(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_453), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_446)
    );

CNN_Single_Layer    single_454(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_454), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_445)
    );

CNN_Single_Layer    single_455(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_455), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_444)
    );

CNN_Single_Layer    single_456(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_456), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_443)
    );

CNN_Single_Layer    single_457(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_457), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_442)
    );

CNN_Single_Layer    single_458(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_458), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_441)
    );

CNN_Single_Layer    single_459(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_459), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_440)
    );

CNN_Single_Layer    single_460(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_460), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_439)
    );

CNN_Single_Layer    single_461(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_461), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_438)
    );

CNN_Single_Layer    single_462(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_462), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_437)
    );

CNN_Single_Layer    single_463(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_463), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_436)
    );

CNN_Single_Layer    single_464(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_464), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_435)
    );

CNN_Single_Layer    single_465(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_465), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_434)
    );

CNN_Single_Layer    single_466(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_466), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_433)
    );

CNN_Single_Layer    single_467(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_467), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_432)
    );

CNN_Single_Layer    single_468(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_468), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_431)
    );

CNN_Single_Layer    single_469(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_469), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_430)
    );

CNN_Single_Layer    single_470(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_470), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_429)
    );

CNN_Single_Layer    single_471(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_471), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_428)
    );

CNN_Single_Layer    single_472(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_472), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_427)
    );

CNN_Single_Layer    single_473(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_473), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_426)
    );

CNN_Single_Layer    single_474(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_474), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_425)
    );

CNN_Single_Layer    single_475(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_475), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_424)
    );

CNN_Single_Layer    single_476(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_476), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_423)
    );

CNN_Single_Layer    single_477(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_477), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_422)
    );

CNN_Single_Layer    single_478(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_478), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_421)
    );

CNN_Single_Layer    single_479(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_479), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_420)
    );

CNN_Single_Layer    single_480(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_480), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_419)
    );

CNN_Single_Layer    single_481(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_481), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_418)
    );

CNN_Single_Layer    single_482(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_482), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_417)
    );

CNN_Single_Layer    single_483(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_483), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_416)
    );

CNN_Single_Layer    single_484(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_484), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_415)
    );

CNN_Single_Layer    single_485(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_485), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_414)
    );

CNN_Single_Layer    single_486(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_486), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_413)
    );

CNN_Single_Layer    single_487(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_487), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_412)
    );

CNN_Single_Layer    single_488(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_488), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_411)
    );

CNN_Single_Layer    single_489(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_489), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_410)
    );

CNN_Single_Layer    single_490(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_490), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_409)
    );

CNN_Single_Layer    single_491(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_491), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_408)
    );

CNN_Single_Layer    single_492(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_492), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_407)
    );

CNN_Single_Layer    single_493(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_493), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_406)
    );

CNN_Single_Layer    single_494(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_494), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_405)
    );

CNN_Single_Layer    single_495(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_495), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_404)
    );

CNN_Single_Layer    single_496(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_496), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_403)
    );

CNN_Single_Layer    single_497(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_497), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_402)
    );

CNN_Single_Layer    single_498(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_498), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_401)
    );

CNN_Single_Layer    single_499(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_499), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_400)
    );

CNN_Single_Layer    single_500(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_500), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_399)
    );

CNN_Single_Layer    single_501(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_501), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_398)
    );

CNN_Single_Layer    single_502(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_502), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_397)
    );

CNN_Single_Layer    single_503(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_503), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_396)
    );

CNN_Single_Layer    single_504(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_504), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_395)
    );

CNN_Single_Layer    single_505(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_505), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_394)
    );

CNN_Single_Layer    single_506(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_506), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_393)
    );

CNN_Single_Layer    single_507(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_507), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_392)
    );

CNN_Single_Layer    single_508(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_508), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_391)
    );

CNN_Single_Layer    single_509(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_509), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_390)
    );

CNN_Single_Layer    single_510(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_510), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_389)
    );

CNN_Single_Layer    single_511(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_511), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_388)
    );

CNN_Single_Layer    single_512(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_512), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_387)
    );

CNN_Single_Layer    single_513(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_513), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_386)
    );

CNN_Single_Layer    single_514(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_514), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_385)
    );

CNN_Single_Layer    single_515(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_515), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_384)
    );

CNN_Single_Layer    single_516(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_516), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_383)
    );

CNN_Single_Layer    single_517(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_517), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_382)
    );

CNN_Single_Layer    single_518(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_518), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_381)
    );

CNN_Single_Layer    single_519(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_519), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_380)
    );

CNN_Single_Layer    single_520(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_520), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_379)
    );

CNN_Single_Layer    single_521(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_521), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_378)
    );

CNN_Single_Layer    single_522(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_522), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_377)
    );

CNN_Single_Layer    single_523(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_523), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_376)
    );

CNN_Single_Layer    single_524(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_524), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_375)
    );

CNN_Single_Layer    single_525(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_525), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_374)
    );

CNN_Single_Layer    single_526(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_526), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_373)
    );

CNN_Single_Layer    single_527(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_527), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_372)
    );

CNN_Single_Layer    single_528(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_528), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_371)
    );

CNN_Single_Layer    single_529(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_529), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_370)
    );

CNN_Single_Layer    single_530(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_530), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_369)
    );

CNN_Single_Layer    single_531(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_531), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_368)
    );

CNN_Single_Layer    single_532(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_532), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_367)
    );

CNN_Single_Layer    single_533(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_533), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_366)
    );

CNN_Single_Layer    single_534(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_534), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_365)
    );

CNN_Single_Layer    single_535(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_535), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_364)
    );

CNN_Single_Layer    single_536(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_536), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_363)
    );

CNN_Single_Layer    single_537(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_537), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_362)
    );

CNN_Single_Layer    single_538(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_538), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_361)
    );

CNN_Single_Layer    single_539(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_539), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_360)
    );

CNN_Single_Layer    single_540(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_540), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_359)
    );

CNN_Single_Layer    single_541(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_541), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_358)
    );

CNN_Single_Layer    single_542(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_542), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_357)
    );

CNN_Single_Layer    single_543(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_543), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_356)
    );

CNN_Single_Layer    single_544(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_544), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_355)
    );

CNN_Single_Layer    single_545(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_545), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_354)
    );

CNN_Single_Layer    single_546(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_546), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_353)
    );

CNN_Single_Layer    single_547(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_547), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_352)
    );

CNN_Single_Layer    single_548(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_548), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_351)
    );

CNN_Single_Layer    single_549(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_549), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_350)
    );

CNN_Single_Layer    single_550(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_550), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_349)
    );

CNN_Single_Layer    single_551(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_551), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_348)
    );

CNN_Single_Layer    single_552(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_552), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_347)
    );

CNN_Single_Layer    single_553(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_553), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_346)
    );

CNN_Single_Layer    single_554(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_554), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_345)
    );

CNN_Single_Layer    single_555(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_555), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_344)
    );

CNN_Single_Layer    single_556(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_556), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_343)
    );

CNN_Single_Layer    single_557(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_557), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_342)
    );

CNN_Single_Layer    single_558(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_558), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_341)
    );

CNN_Single_Layer    single_559(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_559), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_340)
    );

CNN_Single_Layer    single_560(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_560), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_339)
    );

CNN_Single_Layer    single_561(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_561), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_338)
    );

CNN_Single_Layer    single_562(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_562), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_337)
    );

CNN_Single_Layer    single_563(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_563), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_336)
    );

CNN_Single_Layer    single_564(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_564), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_335)
    );

CNN_Single_Layer    single_565(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_565), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_334)
    );

CNN_Single_Layer    single_566(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_566), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_333)
    );

CNN_Single_Layer    single_567(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_567), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_332)
    );

CNN_Single_Layer    single_568(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_568), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_331)
    );

CNN_Single_Layer    single_569(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_569), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_330)
    );

CNN_Single_Layer    single_570(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_570), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_329)
    );

CNN_Single_Layer    single_571(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_571), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_328)
    );

CNN_Single_Layer    single_572(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_572), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_327)
    );

CNN_Single_Layer    single_573(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_573), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_326)
    );

CNN_Single_Layer    single_574(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_574), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_325)
    );

CNN_Single_Layer    single_575(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_575), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_324)
    );

CNN_Single_Layer    single_576(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_576), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_323)
    );

CNN_Single_Layer    single_577(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_577), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_322)
    );

CNN_Single_Layer    single_578(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_578), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_321)
    );

CNN_Single_Layer    single_579(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_579), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_320)
    );

CNN_Single_Layer    single_580(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_580), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_319)
    );

CNN_Single_Layer    single_581(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_581), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_318)
    );

CNN_Single_Layer    single_582(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_582), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_317)
    );

CNN_Single_Layer    single_583(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_583), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_316)
    );

CNN_Single_Layer    single_584(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_584), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_315)
    );

CNN_Single_Layer    single_585(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_585), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_314)
    );

CNN_Single_Layer    single_586(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_586), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_313)
    );

CNN_Single_Layer    single_587(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_587), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_312)
    );

CNN_Single_Layer    single_588(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_588), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_311)
    );

CNN_Single_Layer    single_589(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_589), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_310)
    );

CNN_Single_Layer    single_590(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_590), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_309)
    );

CNN_Single_Layer    single_591(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_591), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_308)
    );

CNN_Single_Layer    single_592(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_592), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_307)
    );

CNN_Single_Layer    single_593(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_593), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_306)
    );

CNN_Single_Layer    single_594(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_594), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_305)
    );

CNN_Single_Layer    single_595(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_595), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_304)
    );

CNN_Single_Layer    single_596(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_596), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_303)
    );

CNN_Single_Layer    single_597(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_597), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_302)
    );

CNN_Single_Layer    single_598(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_598), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_301)
    );

CNN_Single_Layer    single_599(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_599), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_300)
    );

CNN_Single_Layer    single_600(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_600), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_299)
    );

CNN_Single_Layer    single_601(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_601), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_298)
    );

CNN_Single_Layer    single_602(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_602), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_297)
    );

CNN_Single_Layer    single_603(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_603), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_296)
    );

CNN_Single_Layer    single_604(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_604), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_295)
    );

CNN_Single_Layer    single_605(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_605), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_294)
    );

CNN_Single_Layer    single_606(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_606), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_293)
    );

CNN_Single_Layer    single_607(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_607), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_292)
    );

CNN_Single_Layer    single_608(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_608), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_291)
    );

CNN_Single_Layer    single_609(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_609), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_290)
    );

CNN_Single_Layer    single_610(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_610), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_289)
    );

CNN_Single_Layer    single_611(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_611), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_288)
    );

CNN_Single_Layer    single_612(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_612), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_287)
    );

CNN_Single_Layer    single_613(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_613), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_286)
    );

CNN_Single_Layer    single_614(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_614), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_285)
    );

CNN_Single_Layer    single_615(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_615), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_284)
    );

CNN_Single_Layer    single_616(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_616), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_283)
    );

CNN_Single_Layer    single_617(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_617), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_282)
    );

CNN_Single_Layer    single_618(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_618), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_281)
    );

CNN_Single_Layer    single_619(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_619), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_280)
    );

CNN_Single_Layer    single_620(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_620), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_279)
    );

CNN_Single_Layer    single_621(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_621), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_278)
    );

CNN_Single_Layer    single_622(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_622), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_277)
    );

CNN_Single_Layer    single_623(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_623), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_276)
    );

CNN_Single_Layer    single_624(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_624), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_275)
    );

CNN_Single_Layer    single_625(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_625), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_274)
    );

CNN_Single_Layer    single_626(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_626), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_273)
    );

CNN_Single_Layer    single_627(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_627), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_272)
    );

CNN_Single_Layer    single_628(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_628), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_271)
    );

CNN_Single_Layer    single_629(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_629), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_270)
    );

CNN_Single_Layer    single_630(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_630), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_269)
    );

CNN_Single_Layer    single_631(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_631), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_268)
    );

CNN_Single_Layer    single_632(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_632), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_267)
    );

CNN_Single_Layer    single_633(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_633), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_266)
    );

CNN_Single_Layer    single_634(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_634), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_265)
    );

CNN_Single_Layer    single_635(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_635), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_264)
    );

CNN_Single_Layer    single_636(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_636), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_263)
    );

CNN_Single_Layer    single_637(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_637), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_262)
    );

CNN_Single_Layer    single_638(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_638), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_261)
    );

CNN_Single_Layer    single_639(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_639), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_260)
    );

CNN_Single_Layer    single_640(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_640), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_259)
    );

CNN_Single_Layer    single_641(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_641), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_258)
    );

CNN_Single_Layer    single_642(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_642), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_257)
    );

CNN_Single_Layer    single_643(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_643), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_256)
    );

CNN_Single_Layer    single_644(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_644), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_255)
    );

CNN_Single_Layer    single_645(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_645), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_254)
    );

CNN_Single_Layer    single_646(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_646), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_253)
    );

CNN_Single_Layer    single_647(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_647), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_252)
    );

CNN_Single_Layer    single_648(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_648), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_251)
    );

CNN_Single_Layer    single_649(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_649), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_250)
    );

CNN_Single_Layer    single_650(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_650), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_249)
    );

CNN_Single_Layer    single_651(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_651), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_248)
    );

CNN_Single_Layer    single_652(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_652), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_247)
    );

CNN_Single_Layer    single_653(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_653), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_246)
    );

CNN_Single_Layer    single_654(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_654), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_245)
    );

CNN_Single_Layer    single_655(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_655), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_244)
    );

CNN_Single_Layer    single_656(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_656), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_243)
    );

CNN_Single_Layer    single_657(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_657), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_242)
    );

CNN_Single_Layer    single_658(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_658), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_241)
    );

CNN_Single_Layer    single_659(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_659), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_240)
    );

CNN_Single_Layer    single_660(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_660), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_239)
    );

CNN_Single_Layer    single_661(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_661), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_238)
    );

CNN_Single_Layer    single_662(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_662), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_237)
    );

CNN_Single_Layer    single_663(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_663), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_236)
    );

CNN_Single_Layer    single_664(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_664), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_235)
    );

CNN_Single_Layer    single_665(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_665), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_234)
    );

CNN_Single_Layer    single_666(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_666), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_233)
    );

CNN_Single_Layer    single_667(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_667), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_232)
    );

CNN_Single_Layer    single_668(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_668), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_231)
    );

CNN_Single_Layer    single_669(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_669), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_230)
    );

CNN_Single_Layer    single_670(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_670), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_229)
    );

CNN_Single_Layer    single_671(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_671), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_228)
    );

CNN_Single_Layer    single_672(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_672), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_227)
    );

CNN_Single_Layer    single_673(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_673), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_226)
    );

CNN_Single_Layer    single_674(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_674), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_225)
    );

CNN_Single_Layer    single_675(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_675), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_224)
    );

CNN_Single_Layer    single_676(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_676), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_223)
    );

CNN_Single_Layer    single_677(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_677), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_222)
    );

CNN_Single_Layer    single_678(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_678), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_221)
    );

CNN_Single_Layer    single_679(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_679), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_220)
    );

CNN_Single_Layer    single_680(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_680), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_219)
    );

CNN_Single_Layer    single_681(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_681), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_218)
    );

CNN_Single_Layer    single_682(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_682), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_217)
    );

CNN_Single_Layer    single_683(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_683), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_216)
    );

CNN_Single_Layer    single_684(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_684), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_215)
    );

CNN_Single_Layer    single_685(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_685), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_214)
    );

CNN_Single_Layer    single_686(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_686), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_213)
    );

CNN_Single_Layer    single_687(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_687), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_212)
    );

CNN_Single_Layer    single_688(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_688), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_211)
    );

CNN_Single_Layer    single_689(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_689), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_210)
    );

CNN_Single_Layer    single_690(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_690), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_209)
    );

CNN_Single_Layer    single_691(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_691), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_208)
    );

CNN_Single_Layer    single_692(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_692), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_207)
    );

CNN_Single_Layer    single_693(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_693), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_206)
    );

CNN_Single_Layer    single_694(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_694), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_205)
    );

CNN_Single_Layer    single_695(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_695), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_204)
    );

CNN_Single_Layer    single_696(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_696), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_203)
    );

CNN_Single_Layer    single_697(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_697), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_202)
    );

CNN_Single_Layer    single_698(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_698), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_201)
    );

CNN_Single_Layer    single_699(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_699), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_200)
    );

CNN_Single_Layer    single_700(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_700), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_199)
    );

CNN_Single_Layer    single_701(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_701), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_198)
    );

CNN_Single_Layer    single_702(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_702), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_197)
    );

CNN_Single_Layer    single_703(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_703), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_196)
    );

CNN_Single_Layer    single_704(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_704), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_195)
    );

CNN_Single_Layer    single_705(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_705), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_194)
    );

CNN_Single_Layer    single_706(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_706), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_193)
    );

CNN_Single_Layer    single_707(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_707), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_192)
    );

CNN_Single_Layer    single_708(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_708), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_191)
    );

CNN_Single_Layer    single_709(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_709), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_190)
    );

CNN_Single_Layer    single_710(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_710), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_189)
    );

CNN_Single_Layer    single_711(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_711), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_188)
    );

CNN_Single_Layer    single_712(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_712), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_187)
    );

CNN_Single_Layer    single_713(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_713), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_186)
    );

CNN_Single_Layer    single_714(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_714), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_185)
    );

CNN_Single_Layer    single_715(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_715), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_184)
    );

CNN_Single_Layer    single_716(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_716), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_183)
    );

CNN_Single_Layer    single_717(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_717), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_182)
    );

CNN_Single_Layer    single_718(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_718), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_181)
    );

CNN_Single_Layer    single_719(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_719), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_180)
    );

CNN_Single_Layer    single_720(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_720), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_179)
    );

CNN_Single_Layer    single_721(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_721), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_178)
    );

CNN_Single_Layer    single_722(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_722), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_177)
    );

CNN_Single_Layer    single_723(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_723), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_176)
    );

CNN_Single_Layer    single_724(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_724), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_175)
    );

CNN_Single_Layer    single_725(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_725), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_174)
    );

CNN_Single_Layer    single_726(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_726), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_173)
    );

CNN_Single_Layer    single_727(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_727), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_172)
    );

CNN_Single_Layer    single_728(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_728), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_171)
    );

CNN_Single_Layer    single_729(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_729), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_170)
    );

CNN_Single_Layer    single_730(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_730), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_169)
    );

CNN_Single_Layer    single_731(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_731), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_168)
    );

CNN_Single_Layer    single_732(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_732), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_167)
    );

CNN_Single_Layer    single_733(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_733), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_166)
    );

CNN_Single_Layer    single_734(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_734), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_165)
    );

CNN_Single_Layer    single_735(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_735), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_164)
    );

CNN_Single_Layer    single_736(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_736), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_163)
    );

CNN_Single_Layer    single_737(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_737), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_162)
    );

CNN_Single_Layer    single_738(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_738), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_161)
    );

CNN_Single_Layer    single_739(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_739), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_160)
    );

CNN_Single_Layer    single_740(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_740), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_159)
    );

CNN_Single_Layer    single_741(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_741), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_158)
    );

CNN_Single_Layer    single_742(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_742), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_157)
    );

CNN_Single_Layer    single_743(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_743), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_156)
    );

CNN_Single_Layer    single_744(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_744), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_155)
    );

CNN_Single_Layer    single_745(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_745), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_154)
    );

CNN_Single_Layer    single_746(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_746), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_153)
    );

CNN_Single_Layer    single_747(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_747), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_152)
    );

CNN_Single_Layer    single_748(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_748), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_151)
    );

CNN_Single_Layer    single_749(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_749), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_150)
    );

CNN_Single_Layer    single_750(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_750), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_149)
    );

CNN_Single_Layer    single_751(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_751), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_148)
    );

CNN_Single_Layer    single_752(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_752), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_147)
    );

CNN_Single_Layer    single_753(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_753), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_146)
    );

CNN_Single_Layer    single_754(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_754), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_145)
    );

CNN_Single_Layer    single_755(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_755), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_144)
    );

CNN_Single_Layer    single_756(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_756), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_143)
    );

CNN_Single_Layer    single_757(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_757), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_142)
    );

CNN_Single_Layer    single_758(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_758), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_141)
    );

CNN_Single_Layer    single_759(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_759), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_140)
    );

CNN_Single_Layer    single_760(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_760), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_139)
    );

CNN_Single_Layer    single_761(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_761), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_138)
    );

CNN_Single_Layer    single_762(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_762), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_137)
    );

CNN_Single_Layer    single_763(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_763), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_136)
    );

CNN_Single_Layer    single_764(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_764), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_135)
    );

CNN_Single_Layer    single_765(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_765), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_134)
    );

CNN_Single_Layer    single_766(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_766), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_133)
    );

CNN_Single_Layer    single_767(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_767), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_132)
    );

CNN_Single_Layer    single_768(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_768), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_131)
    );

CNN_Single_Layer    single_769(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_769), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_130)
    );

CNN_Single_Layer    single_770(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_770), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_129)
    );

CNN_Single_Layer    single_771(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_771), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_128)
    );

CNN_Single_Layer    single_772(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_772), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_127)
    );

CNN_Single_Layer    single_773(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_773), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_126)
    );

CNN_Single_Layer    single_774(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_774), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_125)
    );

CNN_Single_Layer    single_775(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_775), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_124)
    );

CNN_Single_Layer    single_776(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_776), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_123)
    );

CNN_Single_Layer    single_777(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_777), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_122)
    );

CNN_Single_Layer    single_778(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_778), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_121)
    );

CNN_Single_Layer    single_779(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_779), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_120)
    );

CNN_Single_Layer    single_780(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_780), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_119)
    );

CNN_Single_Layer    single_781(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_781), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_118)
    );

CNN_Single_Layer    single_782(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_782), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_117)
    );

CNN_Single_Layer    single_783(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_783), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_116)
    );

CNN_Single_Layer    single_784(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_784), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_115)
    );

CNN_Single_Layer    single_785(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_785), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_114)
    );

CNN_Single_Layer    single_786(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_786), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_113)
    );

CNN_Single_Layer    single_787(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_787), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_112)
    );

CNN_Single_Layer    single_788(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_788), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_111)
    );

CNN_Single_Layer    single_789(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_789), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_110)
    );

CNN_Single_Layer    single_790(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_790), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_109)
    );

CNN_Single_Layer    single_791(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_791), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_108)
    );

CNN_Single_Layer    single_792(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_792), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_107)
    );

CNN_Single_Layer    single_793(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_793), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_106)
    );

CNN_Single_Layer    single_794(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_794), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_105)
    );

CNN_Single_Layer    single_795(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_795), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_104)
    );

CNN_Single_Layer    single_796(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_796), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_103)
    );

CNN_Single_Layer    single_797(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_797), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_102)
    );

CNN_Single_Layer    single_798(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_798), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_101)
    );

CNN_Single_Layer    single_799(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_799), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_100)
    );

CNN_Single_Layer    single_800(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_800), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_99)
    );

CNN_Single_Layer    single_801(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_801), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_98)
    );

CNN_Single_Layer    single_802(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_802), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_97)
    );

CNN_Single_Layer    single_803(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_803), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_96)
    );

CNN_Single_Layer    single_804(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_804), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_95)
    );

CNN_Single_Layer    single_805(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_805), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_94)
    );

CNN_Single_Layer    single_806(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_806), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_93)
    );

CNN_Single_Layer    single_807(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_807), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_92)
    );

CNN_Single_Layer    single_808(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_808), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_91)
    );

CNN_Single_Layer    single_809(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_809), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_90)
    );

CNN_Single_Layer    single_810(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_810), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_89)
    );

CNN_Single_Layer    single_811(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_811), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_88)
    );

CNN_Single_Layer    single_812(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_812), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_87)
    );

CNN_Single_Layer    single_813(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_813), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_86)
    );

CNN_Single_Layer    single_814(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_814), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_85)
    );

CNN_Single_Layer    single_815(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_815), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_84)
    );

CNN_Single_Layer    single_816(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_816), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_83)
    );

CNN_Single_Layer    single_817(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_817), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_82)
    );

CNN_Single_Layer    single_818(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_818), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_81)
    );

CNN_Single_Layer    single_819(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_819), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_80)
    );

CNN_Single_Layer    single_820(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_820), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_79)
    );

CNN_Single_Layer    single_821(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_821), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_78)
    );

CNN_Single_Layer    single_822(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_822), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_77)
    );

CNN_Single_Layer    single_823(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_823), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_76)
    );

CNN_Single_Layer    single_824(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_824), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_75)
    );

CNN_Single_Layer    single_825(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_825), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_74)
    );

CNN_Single_Layer    single_826(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_826), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_73)
    );

CNN_Single_Layer    single_827(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_827), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_72)
    );

CNN_Single_Layer    single_828(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_828), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_71)
    );

CNN_Single_Layer    single_829(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_829), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_70)
    );

CNN_Single_Layer    single_830(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_830), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_69)
    );

CNN_Single_Layer    single_831(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_831), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_68)
    );

CNN_Single_Layer    single_832(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_832), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_67)
    );

CNN_Single_Layer    single_833(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_833), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_66)
    );

CNN_Single_Layer    single_834(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_834), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_65)
    );

CNN_Single_Layer    single_835(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_835), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_64)
    );

CNN_Single_Layer    single_836(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_836), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_63)
    );

CNN_Single_Layer    single_837(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_837), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_62)
    );

CNN_Single_Layer    single_838(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_838), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_61)
    );

CNN_Single_Layer    single_839(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_839), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_60)
    );

CNN_Single_Layer    single_840(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_840), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_59)
    );

CNN_Single_Layer    single_841(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_841), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_58)
    );

CNN_Single_Layer    single_842(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_842), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_57)
    );

CNN_Single_Layer    single_843(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_843), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_56)
    );

CNN_Single_Layer    single_844(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_844), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_55)
    );

CNN_Single_Layer    single_845(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_845), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_54)
    );

CNN_Single_Layer    single_846(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_846), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_53)
    );

CNN_Single_Layer    single_847(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_847), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_52)
    );

CNN_Single_Layer    single_848(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_848), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_51)
    );

CNN_Single_Layer    single_849(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_849), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_50)
    );

CNN_Single_Layer    single_850(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_850), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_49)
    );

CNN_Single_Layer    single_851(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_851), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_48)
    );

CNN_Single_Layer    single_852(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_852), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_47)
    );

CNN_Single_Layer    single_853(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_853), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_46)
    );

CNN_Single_Layer    single_854(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_854), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_45)
    );

CNN_Single_Layer    single_855(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_855), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_44)
    );

CNN_Single_Layer    single_856(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_856), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_43)
    );

CNN_Single_Layer    single_857(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_857), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_42)
    );

CNN_Single_Layer    single_858(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_858), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_41)
    );

CNN_Single_Layer    single_859(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_859), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_40)
    );

CNN_Single_Layer    single_860(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_860), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_39)
    );

CNN_Single_Layer    single_861(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_861), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_38)
    );

CNN_Single_Layer    single_862(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_862), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_37)
    );

CNN_Single_Layer    single_863(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_863), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_36)
    );

CNN_Single_Layer    single_864(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_864), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_35)
    );

CNN_Single_Layer    single_865(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_865), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_34)
    );

CNN_Single_Layer    single_866(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_866), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_33)
    );

CNN_Single_Layer    single_867(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_867), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_32)
    );

CNN_Single_Layer    single_868(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_868), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_31)
    );

CNN_Single_Layer    single_869(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_869), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_30)
    );

CNN_Single_Layer    single_870(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_870), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_29)
    );

CNN_Single_Layer    single_871(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_871), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_28)
    );

CNN_Single_Layer    single_872(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_872), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_27)
    );

CNN_Single_Layer    single_873(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_873), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_26)
    );

CNN_Single_Layer    single_874(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_874), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_25)
    );

CNN_Single_Layer    single_875(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_875), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_24)
    );

CNN_Single_Layer    single_876(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_876), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_23)
    );

CNN_Single_Layer    single_877(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_877), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_22)
    );

CNN_Single_Layer    single_878(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_878), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_21)
    );

CNN_Single_Layer    single_879(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_879), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_20)
    );

CNN_Single_Layer    single_880(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_880), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_19)
    );

CNN_Single_Layer    single_881(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_881), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_18)
    );

CNN_Single_Layer    single_882(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_882), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_17)
    );

CNN_Single_Layer    single_883(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_883), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_16)
    );

CNN_Single_Layer    single_884(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_884), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_15)
    );

CNN_Single_Layer    single_885(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_885), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_14)
    );

CNN_Single_Layer    single_886(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_886), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_13)
    );

CNN_Single_Layer    single_887(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_887), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_12)
    );

CNN_Single_Layer    single_888(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_888), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_11)
    );

CNN_Single_Layer    single_889(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_889), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_10)
    );

CNN_Single_Layer    single_890(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_890), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_9)
    );

CNN_Single_Layer    single_891(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_891), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_8)
    );

CNN_Single_Layer    single_892(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_892), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_7)
    );

CNN_Single_Layer    single_893(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_893), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_6)
    );

CNN_Single_Layer    single_894(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_894), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_5)
    );

CNN_Single_Layer    single_895(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_895), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_4)
    );

CNN_Single_Layer    single_896(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_896), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_3)
    );

CNN_Single_Layer    single_897(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_897), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_2)
    );

CNN_Single_Layer    single_898(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_898), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_1)
    );

CNN_Single_Layer    single_899(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_0_899), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_0_0)
    );

always @(*) begin
    Conv_out[0]   <= conv_out_0_0;

    Conv_out[1]   <= conv_out_0_1;

    Conv_out[2]   <= conv_out_0_2;

    Conv_out[3]   <= conv_out_0_3;

    Conv_out[4]   <= conv_out_0_4;

    Conv_out[5]   <= conv_out_0_5;

    Conv_out[6]   <= conv_out_0_6;

    Conv_out[7]   <= conv_out_0_7;

    Conv_out[8]   <= conv_out_0_8;

    Conv_out[9]   <= conv_out_0_9;

    Conv_out[10]   <= conv_out_0_10;

    Conv_out[11]   <= conv_out_0_11;

    Conv_out[12]   <= conv_out_0_12;

    Conv_out[13]   <= conv_out_0_13;

    Conv_out[14]   <= conv_out_0_14;

    Conv_out[15]   <= conv_out_0_15;

    Conv_out[16]   <= conv_out_0_16;

    Conv_out[17]   <= conv_out_0_17;

    Conv_out[18]   <= conv_out_0_18;

    Conv_out[19]   <= conv_out_0_19;

    Conv_out[20]   <= conv_out_0_20;

    Conv_out[21]   <= conv_out_0_21;

    Conv_out[22]   <= conv_out_0_22;

    Conv_out[23]   <= conv_out_0_23;

    Conv_out[24]   <= conv_out_0_24;

    Conv_out[25]   <= conv_out_0_25;

    Conv_out[26]   <= conv_out_0_26;

    Conv_out[27]   <= conv_out_0_27;

    Conv_out[28]   <= conv_out_0_28;

    Conv_out[29]   <= conv_out_0_29;

    Conv_out[30]   <= conv_out_0_30;

    Conv_out[31]   <= conv_out_0_31;

    Conv_out[32]   <= conv_out_0_32;

    Conv_out[33]   <= conv_out_0_33;

    Conv_out[34]   <= conv_out_0_34;

    Conv_out[35]   <= conv_out_0_35;

    Conv_out[36]   <= conv_out_0_36;

    Conv_out[37]   <= conv_out_0_37;

    Conv_out[38]   <= conv_out_0_38;

    Conv_out[39]   <= conv_out_0_39;

    Conv_out[40]   <= conv_out_0_40;

    Conv_out[41]   <= conv_out_0_41;

    Conv_out[42]   <= conv_out_0_42;

    Conv_out[43]   <= conv_out_0_43;

    Conv_out[44]   <= conv_out_0_44;

    Conv_out[45]   <= conv_out_0_45;

    Conv_out[46]   <= conv_out_0_46;

    Conv_out[47]   <= conv_out_0_47;

    Conv_out[48]   <= conv_out_0_48;

    Conv_out[49]   <= conv_out_0_49;

    Conv_out[50]   <= conv_out_0_50;

    Conv_out[51]   <= conv_out_0_51;

    Conv_out[52]   <= conv_out_0_52;

    Conv_out[53]   <= conv_out_0_53;

    Conv_out[54]   <= conv_out_0_54;

    Conv_out[55]   <= conv_out_0_55;

    Conv_out[56]   <= conv_out_0_56;

    Conv_out[57]   <= conv_out_0_57;

    Conv_out[58]   <= conv_out_0_58;

    Conv_out[59]   <= conv_out_0_59;

    Conv_out[60]   <= conv_out_0_60;

    Conv_out[61]   <= conv_out_0_61;

    Conv_out[62]   <= conv_out_0_62;

    Conv_out[63]   <= conv_out_0_63;

    Conv_out[64]   <= conv_out_0_64;

    Conv_out[65]   <= conv_out_0_65;

    Conv_out[66]   <= conv_out_0_66;

    Conv_out[67]   <= conv_out_0_67;

    Conv_out[68]   <= conv_out_0_68;

    Conv_out[69]   <= conv_out_0_69;

    Conv_out[70]   <= conv_out_0_70;

    Conv_out[71]   <= conv_out_0_71;

    Conv_out[72]   <= conv_out_0_72;

    Conv_out[73]   <= conv_out_0_73;

    Conv_out[74]   <= conv_out_0_74;

    Conv_out[75]   <= conv_out_0_75;

    Conv_out[76]   <= conv_out_0_76;

    Conv_out[77]   <= conv_out_0_77;

    Conv_out[78]   <= conv_out_0_78;

    Conv_out[79]   <= conv_out_0_79;

    Conv_out[80]   <= conv_out_0_80;

    Conv_out[81]   <= conv_out_0_81;

    Conv_out[82]   <= conv_out_0_82;

    Conv_out[83]   <= conv_out_0_83;

    Conv_out[84]   <= conv_out_0_84;

    Conv_out[85]   <= conv_out_0_85;

    Conv_out[86]   <= conv_out_0_86;

    Conv_out[87]   <= conv_out_0_87;

    Conv_out[88]   <= conv_out_0_88;

    Conv_out[89]   <= conv_out_0_89;

    Conv_out[90]   <= conv_out_0_90;

    Conv_out[91]   <= conv_out_0_91;

    Conv_out[92]   <= conv_out_0_92;

    Conv_out[93]   <= conv_out_0_93;

    Conv_out[94]   <= conv_out_0_94;

    Conv_out[95]   <= conv_out_0_95;

    Conv_out[96]   <= conv_out_0_96;

    Conv_out[97]   <= conv_out_0_97;

    Conv_out[98]   <= conv_out_0_98;

    Conv_out[99]   <= conv_out_0_99;

    Conv_out[100]   <= conv_out_0_100;

    Conv_out[101]   <= conv_out_0_101;

    Conv_out[102]   <= conv_out_0_102;

    Conv_out[103]   <= conv_out_0_103;

    Conv_out[104]   <= conv_out_0_104;

    Conv_out[105]   <= conv_out_0_105;

    Conv_out[106]   <= conv_out_0_106;

    Conv_out[107]   <= conv_out_0_107;

    Conv_out[108]   <= conv_out_0_108;

    Conv_out[109]   <= conv_out_0_109;

    Conv_out[110]   <= conv_out_0_110;

    Conv_out[111]   <= conv_out_0_111;

    Conv_out[112]   <= conv_out_0_112;

    Conv_out[113]   <= conv_out_0_113;

    Conv_out[114]   <= conv_out_0_114;

    Conv_out[115]   <= conv_out_0_115;

    Conv_out[116]   <= conv_out_0_116;

    Conv_out[117]   <= conv_out_0_117;

    Conv_out[118]   <= conv_out_0_118;

    Conv_out[119]   <= conv_out_0_119;

    Conv_out[120]   <= conv_out_0_120;

    Conv_out[121]   <= conv_out_0_121;

    Conv_out[122]   <= conv_out_0_122;

    Conv_out[123]   <= conv_out_0_123;

    Conv_out[124]   <= conv_out_0_124;

    Conv_out[125]   <= conv_out_0_125;

    Conv_out[126]   <= conv_out_0_126;

    Conv_out[127]   <= conv_out_0_127;

    Conv_out[128]   <= conv_out_0_128;

    Conv_out[129]   <= conv_out_0_129;

    Conv_out[130]   <= conv_out_0_130;

    Conv_out[131]   <= conv_out_0_131;

    Conv_out[132]   <= conv_out_0_132;

    Conv_out[133]   <= conv_out_0_133;

    Conv_out[134]   <= conv_out_0_134;

    Conv_out[135]   <= conv_out_0_135;

    Conv_out[136]   <= conv_out_0_136;

    Conv_out[137]   <= conv_out_0_137;

    Conv_out[138]   <= conv_out_0_138;

    Conv_out[139]   <= conv_out_0_139;

    Conv_out[140]   <= conv_out_0_140;

    Conv_out[141]   <= conv_out_0_141;

    Conv_out[142]   <= conv_out_0_142;

    Conv_out[143]   <= conv_out_0_143;

    Conv_out[144]   <= conv_out_0_144;

    Conv_out[145]   <= conv_out_0_145;

    Conv_out[146]   <= conv_out_0_146;

    Conv_out[147]   <= conv_out_0_147;

    Conv_out[148]   <= conv_out_0_148;

    Conv_out[149]   <= conv_out_0_149;

    Conv_out[150]   <= conv_out_0_150;

    Conv_out[151]   <= conv_out_0_151;

    Conv_out[152]   <= conv_out_0_152;

    Conv_out[153]   <= conv_out_0_153;

    Conv_out[154]   <= conv_out_0_154;

    Conv_out[155]   <= conv_out_0_155;

    Conv_out[156]   <= conv_out_0_156;

    Conv_out[157]   <= conv_out_0_157;

    Conv_out[158]   <= conv_out_0_158;

    Conv_out[159]   <= conv_out_0_159;

    Conv_out[160]   <= conv_out_0_160;

    Conv_out[161]   <= conv_out_0_161;

    Conv_out[162]   <= conv_out_0_162;

    Conv_out[163]   <= conv_out_0_163;

    Conv_out[164]   <= conv_out_0_164;

    Conv_out[165]   <= conv_out_0_165;

    Conv_out[166]   <= conv_out_0_166;

    Conv_out[167]   <= conv_out_0_167;

    Conv_out[168]   <= conv_out_0_168;

    Conv_out[169]   <= conv_out_0_169;

    Conv_out[170]   <= conv_out_0_170;

    Conv_out[171]   <= conv_out_0_171;

    Conv_out[172]   <= conv_out_0_172;

    Conv_out[173]   <= conv_out_0_173;

    Conv_out[174]   <= conv_out_0_174;

    Conv_out[175]   <= conv_out_0_175;

    Conv_out[176]   <= conv_out_0_176;

    Conv_out[177]   <= conv_out_0_177;

    Conv_out[178]   <= conv_out_0_178;

    Conv_out[179]   <= conv_out_0_179;

    Conv_out[180]   <= conv_out_0_180;

    Conv_out[181]   <= conv_out_0_181;

    Conv_out[182]   <= conv_out_0_182;

    Conv_out[183]   <= conv_out_0_183;

    Conv_out[184]   <= conv_out_0_184;

    Conv_out[185]   <= conv_out_0_185;

    Conv_out[186]   <= conv_out_0_186;

    Conv_out[187]   <= conv_out_0_187;

    Conv_out[188]   <= conv_out_0_188;

    Conv_out[189]   <= conv_out_0_189;

    Conv_out[190]   <= conv_out_0_190;

    Conv_out[191]   <= conv_out_0_191;

    Conv_out[192]   <= conv_out_0_192;

    Conv_out[193]   <= conv_out_0_193;

    Conv_out[194]   <= conv_out_0_194;

    Conv_out[195]   <= conv_out_0_195;

    Conv_out[196]   <= conv_out_0_196;

    Conv_out[197]   <= conv_out_0_197;

    Conv_out[198]   <= conv_out_0_198;

    Conv_out[199]   <= conv_out_0_199;

    Conv_out[200]   <= conv_out_0_200;

    Conv_out[201]   <= conv_out_0_201;

    Conv_out[202]   <= conv_out_0_202;

    Conv_out[203]   <= conv_out_0_203;

    Conv_out[204]   <= conv_out_0_204;

    Conv_out[205]   <= conv_out_0_205;

    Conv_out[206]   <= conv_out_0_206;

    Conv_out[207]   <= conv_out_0_207;

    Conv_out[208]   <= conv_out_0_208;

    Conv_out[209]   <= conv_out_0_209;

    Conv_out[210]   <= conv_out_0_210;

    Conv_out[211]   <= conv_out_0_211;

    Conv_out[212]   <= conv_out_0_212;

    Conv_out[213]   <= conv_out_0_213;

    Conv_out[214]   <= conv_out_0_214;

    Conv_out[215]   <= conv_out_0_215;

    Conv_out[216]   <= conv_out_0_216;

    Conv_out[217]   <= conv_out_0_217;

    Conv_out[218]   <= conv_out_0_218;

    Conv_out[219]   <= conv_out_0_219;

    Conv_out[220]   <= conv_out_0_220;

    Conv_out[221]   <= conv_out_0_221;

    Conv_out[222]   <= conv_out_0_222;

    Conv_out[223]   <= conv_out_0_223;

    Conv_out[224]   <= conv_out_0_224;

    Conv_out[225]   <= conv_out_0_225;

    Conv_out[226]   <= conv_out_0_226;

    Conv_out[227]   <= conv_out_0_227;

    Conv_out[228]   <= conv_out_0_228;

    Conv_out[229]   <= conv_out_0_229;

    Conv_out[230]   <= conv_out_0_230;

    Conv_out[231]   <= conv_out_0_231;

    Conv_out[232]   <= conv_out_0_232;

    Conv_out[233]   <= conv_out_0_233;

    Conv_out[234]   <= conv_out_0_234;

    Conv_out[235]   <= conv_out_0_235;

    Conv_out[236]   <= conv_out_0_236;

    Conv_out[237]   <= conv_out_0_237;

    Conv_out[238]   <= conv_out_0_238;

    Conv_out[239]   <= conv_out_0_239;

    Conv_out[240]   <= conv_out_0_240;

    Conv_out[241]   <= conv_out_0_241;

    Conv_out[242]   <= conv_out_0_242;

    Conv_out[243]   <= conv_out_0_243;

    Conv_out[244]   <= conv_out_0_244;

    Conv_out[245]   <= conv_out_0_245;

    Conv_out[246]   <= conv_out_0_246;

    Conv_out[247]   <= conv_out_0_247;

    Conv_out[248]   <= conv_out_0_248;

    Conv_out[249]   <= conv_out_0_249;

    Conv_out[250]   <= conv_out_0_250;

    Conv_out[251]   <= conv_out_0_251;

    Conv_out[252]   <= conv_out_0_252;

    Conv_out[253]   <= conv_out_0_253;

    Conv_out[254]   <= conv_out_0_254;

    Conv_out[255]   <= conv_out_0_255;

    Conv_out[256]   <= conv_out_0_256;

    Conv_out[257]   <= conv_out_0_257;

    Conv_out[258]   <= conv_out_0_258;

    Conv_out[259]   <= conv_out_0_259;

    Conv_out[260]   <= conv_out_0_260;

    Conv_out[261]   <= conv_out_0_261;

    Conv_out[262]   <= conv_out_0_262;

    Conv_out[263]   <= conv_out_0_263;

    Conv_out[264]   <= conv_out_0_264;

    Conv_out[265]   <= conv_out_0_265;

    Conv_out[266]   <= conv_out_0_266;

    Conv_out[267]   <= conv_out_0_267;

    Conv_out[268]   <= conv_out_0_268;

    Conv_out[269]   <= conv_out_0_269;

    Conv_out[270]   <= conv_out_0_270;

    Conv_out[271]   <= conv_out_0_271;

    Conv_out[272]   <= conv_out_0_272;

    Conv_out[273]   <= conv_out_0_273;

    Conv_out[274]   <= conv_out_0_274;

    Conv_out[275]   <= conv_out_0_275;

    Conv_out[276]   <= conv_out_0_276;

    Conv_out[277]   <= conv_out_0_277;

    Conv_out[278]   <= conv_out_0_278;

    Conv_out[279]   <= conv_out_0_279;

    Conv_out[280]   <= conv_out_0_280;

    Conv_out[281]   <= conv_out_0_281;

    Conv_out[282]   <= conv_out_0_282;

    Conv_out[283]   <= conv_out_0_283;

    Conv_out[284]   <= conv_out_0_284;

    Conv_out[285]   <= conv_out_0_285;

    Conv_out[286]   <= conv_out_0_286;

    Conv_out[287]   <= conv_out_0_287;

    Conv_out[288]   <= conv_out_0_288;

    Conv_out[289]   <= conv_out_0_289;

    Conv_out[290]   <= conv_out_0_290;

    Conv_out[291]   <= conv_out_0_291;

    Conv_out[292]   <= conv_out_0_292;

    Conv_out[293]   <= conv_out_0_293;

    Conv_out[294]   <= conv_out_0_294;

    Conv_out[295]   <= conv_out_0_295;

    Conv_out[296]   <= conv_out_0_296;

    Conv_out[297]   <= conv_out_0_297;

    Conv_out[298]   <= conv_out_0_298;

    Conv_out[299]   <= conv_out_0_299;

    Conv_out[300]   <= conv_out_0_300;

    Conv_out[301]   <= conv_out_0_301;

    Conv_out[302]   <= conv_out_0_302;

    Conv_out[303]   <= conv_out_0_303;

    Conv_out[304]   <= conv_out_0_304;

    Conv_out[305]   <= conv_out_0_305;

    Conv_out[306]   <= conv_out_0_306;

    Conv_out[307]   <= conv_out_0_307;

    Conv_out[308]   <= conv_out_0_308;

    Conv_out[309]   <= conv_out_0_309;

    Conv_out[310]   <= conv_out_0_310;

    Conv_out[311]   <= conv_out_0_311;

    Conv_out[312]   <= conv_out_0_312;

    Conv_out[313]   <= conv_out_0_313;

    Conv_out[314]   <= conv_out_0_314;

    Conv_out[315]   <= conv_out_0_315;

    Conv_out[316]   <= conv_out_0_316;

    Conv_out[317]   <= conv_out_0_317;

    Conv_out[318]   <= conv_out_0_318;

    Conv_out[319]   <= conv_out_0_319;

    Conv_out[320]   <= conv_out_0_320;

    Conv_out[321]   <= conv_out_0_321;

    Conv_out[322]   <= conv_out_0_322;

    Conv_out[323]   <= conv_out_0_323;

    Conv_out[324]   <= conv_out_0_324;

    Conv_out[325]   <= conv_out_0_325;

    Conv_out[326]   <= conv_out_0_326;

    Conv_out[327]   <= conv_out_0_327;

    Conv_out[328]   <= conv_out_0_328;

    Conv_out[329]   <= conv_out_0_329;

    Conv_out[330]   <= conv_out_0_330;

    Conv_out[331]   <= conv_out_0_331;

    Conv_out[332]   <= conv_out_0_332;

    Conv_out[333]   <= conv_out_0_333;

    Conv_out[334]   <= conv_out_0_334;

    Conv_out[335]   <= conv_out_0_335;

    Conv_out[336]   <= conv_out_0_336;

    Conv_out[337]   <= conv_out_0_337;

    Conv_out[338]   <= conv_out_0_338;

    Conv_out[339]   <= conv_out_0_339;

    Conv_out[340]   <= conv_out_0_340;

    Conv_out[341]   <= conv_out_0_341;

    Conv_out[342]   <= conv_out_0_342;

    Conv_out[343]   <= conv_out_0_343;

    Conv_out[344]   <= conv_out_0_344;

    Conv_out[345]   <= conv_out_0_345;

    Conv_out[346]   <= conv_out_0_346;

    Conv_out[347]   <= conv_out_0_347;

    Conv_out[348]   <= conv_out_0_348;

    Conv_out[349]   <= conv_out_0_349;

    Conv_out[350]   <= conv_out_0_350;

    Conv_out[351]   <= conv_out_0_351;

    Conv_out[352]   <= conv_out_0_352;

    Conv_out[353]   <= conv_out_0_353;

    Conv_out[354]   <= conv_out_0_354;

    Conv_out[355]   <= conv_out_0_355;

    Conv_out[356]   <= conv_out_0_356;

    Conv_out[357]   <= conv_out_0_357;

    Conv_out[358]   <= conv_out_0_358;

    Conv_out[359]   <= conv_out_0_359;

    Conv_out[360]   <= conv_out_0_360;

    Conv_out[361]   <= conv_out_0_361;

    Conv_out[362]   <= conv_out_0_362;

    Conv_out[363]   <= conv_out_0_363;

    Conv_out[364]   <= conv_out_0_364;

    Conv_out[365]   <= conv_out_0_365;

    Conv_out[366]   <= conv_out_0_366;

    Conv_out[367]   <= conv_out_0_367;

    Conv_out[368]   <= conv_out_0_368;

    Conv_out[369]   <= conv_out_0_369;

    Conv_out[370]   <= conv_out_0_370;

    Conv_out[371]   <= conv_out_0_371;

    Conv_out[372]   <= conv_out_0_372;

    Conv_out[373]   <= conv_out_0_373;

    Conv_out[374]   <= conv_out_0_374;

    Conv_out[375]   <= conv_out_0_375;

    Conv_out[376]   <= conv_out_0_376;

    Conv_out[377]   <= conv_out_0_377;

    Conv_out[378]   <= conv_out_0_378;

    Conv_out[379]   <= conv_out_0_379;

    Conv_out[380]   <= conv_out_0_380;

    Conv_out[381]   <= conv_out_0_381;

    Conv_out[382]   <= conv_out_0_382;

    Conv_out[383]   <= conv_out_0_383;

    Conv_out[384]   <= conv_out_0_384;

    Conv_out[385]   <= conv_out_0_385;

    Conv_out[386]   <= conv_out_0_386;

    Conv_out[387]   <= conv_out_0_387;

    Conv_out[388]   <= conv_out_0_388;

    Conv_out[389]   <= conv_out_0_389;

    Conv_out[390]   <= conv_out_0_390;

    Conv_out[391]   <= conv_out_0_391;

    Conv_out[392]   <= conv_out_0_392;

    Conv_out[393]   <= conv_out_0_393;

    Conv_out[394]   <= conv_out_0_394;

    Conv_out[395]   <= conv_out_0_395;

    Conv_out[396]   <= conv_out_0_396;

    Conv_out[397]   <= conv_out_0_397;

    Conv_out[398]   <= conv_out_0_398;

    Conv_out[399]   <= conv_out_0_399;

    Conv_out[400]   <= conv_out_0_400;

    Conv_out[401]   <= conv_out_0_401;

    Conv_out[402]   <= conv_out_0_402;

    Conv_out[403]   <= conv_out_0_403;

    Conv_out[404]   <= conv_out_0_404;

    Conv_out[405]   <= conv_out_0_405;

    Conv_out[406]   <= conv_out_0_406;

    Conv_out[407]   <= conv_out_0_407;

    Conv_out[408]   <= conv_out_0_408;

    Conv_out[409]   <= conv_out_0_409;

    Conv_out[410]   <= conv_out_0_410;

    Conv_out[411]   <= conv_out_0_411;

    Conv_out[412]   <= conv_out_0_412;

    Conv_out[413]   <= conv_out_0_413;

    Conv_out[414]   <= conv_out_0_414;

    Conv_out[415]   <= conv_out_0_415;

    Conv_out[416]   <= conv_out_0_416;

    Conv_out[417]   <= conv_out_0_417;

    Conv_out[418]   <= conv_out_0_418;

    Conv_out[419]   <= conv_out_0_419;

    Conv_out[420]   <= conv_out_0_420;

    Conv_out[421]   <= conv_out_0_421;

    Conv_out[422]   <= conv_out_0_422;

    Conv_out[423]   <= conv_out_0_423;

    Conv_out[424]   <= conv_out_0_424;

    Conv_out[425]   <= conv_out_0_425;

    Conv_out[426]   <= conv_out_0_426;

    Conv_out[427]   <= conv_out_0_427;

    Conv_out[428]   <= conv_out_0_428;

    Conv_out[429]   <= conv_out_0_429;

    Conv_out[430]   <= conv_out_0_430;

    Conv_out[431]   <= conv_out_0_431;

    Conv_out[432]   <= conv_out_0_432;

    Conv_out[433]   <= conv_out_0_433;

    Conv_out[434]   <= conv_out_0_434;

    Conv_out[435]   <= conv_out_0_435;

    Conv_out[436]   <= conv_out_0_436;

    Conv_out[437]   <= conv_out_0_437;

    Conv_out[438]   <= conv_out_0_438;

    Conv_out[439]   <= conv_out_0_439;

    Conv_out[440]   <= conv_out_0_440;

    Conv_out[441]   <= conv_out_0_441;

    Conv_out[442]   <= conv_out_0_442;

    Conv_out[443]   <= conv_out_0_443;

    Conv_out[444]   <= conv_out_0_444;

    Conv_out[445]   <= conv_out_0_445;

    Conv_out[446]   <= conv_out_0_446;

    Conv_out[447]   <= conv_out_0_447;

    Conv_out[448]   <= conv_out_0_448;

    Conv_out[449]   <= conv_out_0_449;

    Conv_out[450]   <= conv_out_0_450;

    Conv_out[451]   <= conv_out_0_451;

    Conv_out[452]   <= conv_out_0_452;

    Conv_out[453]   <= conv_out_0_453;

    Conv_out[454]   <= conv_out_0_454;

    Conv_out[455]   <= conv_out_0_455;

    Conv_out[456]   <= conv_out_0_456;

    Conv_out[457]   <= conv_out_0_457;

    Conv_out[458]   <= conv_out_0_458;

    Conv_out[459]   <= conv_out_0_459;

    Conv_out[460]   <= conv_out_0_460;

    Conv_out[461]   <= conv_out_0_461;

    Conv_out[462]   <= conv_out_0_462;

    Conv_out[463]   <= conv_out_0_463;

    Conv_out[464]   <= conv_out_0_464;

    Conv_out[465]   <= conv_out_0_465;

    Conv_out[466]   <= conv_out_0_466;

    Conv_out[467]   <= conv_out_0_467;

    Conv_out[468]   <= conv_out_0_468;

    Conv_out[469]   <= conv_out_0_469;

    Conv_out[470]   <= conv_out_0_470;

    Conv_out[471]   <= conv_out_0_471;

    Conv_out[472]   <= conv_out_0_472;

    Conv_out[473]   <= conv_out_0_473;

    Conv_out[474]   <= conv_out_0_474;

    Conv_out[475]   <= conv_out_0_475;

    Conv_out[476]   <= conv_out_0_476;

    Conv_out[477]   <= conv_out_0_477;

    Conv_out[478]   <= conv_out_0_478;

    Conv_out[479]   <= conv_out_0_479;

    Conv_out[480]   <= conv_out_0_480;

    Conv_out[481]   <= conv_out_0_481;

    Conv_out[482]   <= conv_out_0_482;

    Conv_out[483]   <= conv_out_0_483;

    Conv_out[484]   <= conv_out_0_484;

    Conv_out[485]   <= conv_out_0_485;

    Conv_out[486]   <= conv_out_0_486;

    Conv_out[487]   <= conv_out_0_487;

    Conv_out[488]   <= conv_out_0_488;

    Conv_out[489]   <= conv_out_0_489;

    Conv_out[490]   <= conv_out_0_490;

    Conv_out[491]   <= conv_out_0_491;

    Conv_out[492]   <= conv_out_0_492;

    Conv_out[493]   <= conv_out_0_493;

    Conv_out[494]   <= conv_out_0_494;

    Conv_out[495]   <= conv_out_0_495;

    Conv_out[496]   <= conv_out_0_496;

    Conv_out[497]   <= conv_out_0_497;

    Conv_out[498]   <= conv_out_0_498;

    Conv_out[499]   <= conv_out_0_499;

    Conv_out[500]   <= conv_out_0_500;

    Conv_out[501]   <= conv_out_0_501;

    Conv_out[502]   <= conv_out_0_502;

    Conv_out[503]   <= conv_out_0_503;

    Conv_out[504]   <= conv_out_0_504;

    Conv_out[505]   <= conv_out_0_505;

    Conv_out[506]   <= conv_out_0_506;

    Conv_out[507]   <= conv_out_0_507;

    Conv_out[508]   <= conv_out_0_508;

    Conv_out[509]   <= conv_out_0_509;

    Conv_out[510]   <= conv_out_0_510;

    Conv_out[511]   <= conv_out_0_511;

    Conv_out[512]   <= conv_out_0_512;

    Conv_out[513]   <= conv_out_0_513;

    Conv_out[514]   <= conv_out_0_514;

    Conv_out[515]   <= conv_out_0_515;

    Conv_out[516]   <= conv_out_0_516;

    Conv_out[517]   <= conv_out_0_517;

    Conv_out[518]   <= conv_out_0_518;

    Conv_out[519]   <= conv_out_0_519;

    Conv_out[520]   <= conv_out_0_520;

    Conv_out[521]   <= conv_out_0_521;

    Conv_out[522]   <= conv_out_0_522;

    Conv_out[523]   <= conv_out_0_523;

    Conv_out[524]   <= conv_out_0_524;

    Conv_out[525]   <= conv_out_0_525;

    Conv_out[526]   <= conv_out_0_526;

    Conv_out[527]   <= conv_out_0_527;

    Conv_out[528]   <= conv_out_0_528;

    Conv_out[529]   <= conv_out_0_529;

    Conv_out[530]   <= conv_out_0_530;

    Conv_out[531]   <= conv_out_0_531;

    Conv_out[532]   <= conv_out_0_532;

    Conv_out[533]   <= conv_out_0_533;

    Conv_out[534]   <= conv_out_0_534;

    Conv_out[535]   <= conv_out_0_535;

    Conv_out[536]   <= conv_out_0_536;

    Conv_out[537]   <= conv_out_0_537;

    Conv_out[538]   <= conv_out_0_538;

    Conv_out[539]   <= conv_out_0_539;

    Conv_out[540]   <= conv_out_0_540;

    Conv_out[541]   <= conv_out_0_541;

    Conv_out[542]   <= conv_out_0_542;

    Conv_out[543]   <= conv_out_0_543;

    Conv_out[544]   <= conv_out_0_544;

    Conv_out[545]   <= conv_out_0_545;

    Conv_out[546]   <= conv_out_0_546;

    Conv_out[547]   <= conv_out_0_547;

    Conv_out[548]   <= conv_out_0_548;

    Conv_out[549]   <= conv_out_0_549;

    Conv_out[550]   <= conv_out_0_550;

    Conv_out[551]   <= conv_out_0_551;

    Conv_out[552]   <= conv_out_0_552;

    Conv_out[553]   <= conv_out_0_553;

    Conv_out[554]   <= conv_out_0_554;

    Conv_out[555]   <= conv_out_0_555;

    Conv_out[556]   <= conv_out_0_556;

    Conv_out[557]   <= conv_out_0_557;

    Conv_out[558]   <= conv_out_0_558;

    Conv_out[559]   <= conv_out_0_559;

    Conv_out[560]   <= conv_out_0_560;

    Conv_out[561]   <= conv_out_0_561;

    Conv_out[562]   <= conv_out_0_562;

    Conv_out[563]   <= conv_out_0_563;

    Conv_out[564]   <= conv_out_0_564;

    Conv_out[565]   <= conv_out_0_565;

    Conv_out[566]   <= conv_out_0_566;

    Conv_out[567]   <= conv_out_0_567;

    Conv_out[568]   <= conv_out_0_568;

    Conv_out[569]   <= conv_out_0_569;

    Conv_out[570]   <= conv_out_0_570;

    Conv_out[571]   <= conv_out_0_571;

    Conv_out[572]   <= conv_out_0_572;

    Conv_out[573]   <= conv_out_0_573;

    Conv_out[574]   <= conv_out_0_574;

    Conv_out[575]   <= conv_out_0_575;

    Conv_out[576]   <= conv_out_0_576;

    Conv_out[577]   <= conv_out_0_577;

    Conv_out[578]   <= conv_out_0_578;

    Conv_out[579]   <= conv_out_0_579;

    Conv_out[580]   <= conv_out_0_580;

    Conv_out[581]   <= conv_out_0_581;

    Conv_out[582]   <= conv_out_0_582;

    Conv_out[583]   <= conv_out_0_583;

    Conv_out[584]   <= conv_out_0_584;

    Conv_out[585]   <= conv_out_0_585;

    Conv_out[586]   <= conv_out_0_586;

    Conv_out[587]   <= conv_out_0_587;

    Conv_out[588]   <= conv_out_0_588;

    Conv_out[589]   <= conv_out_0_589;

    Conv_out[590]   <= conv_out_0_590;

    Conv_out[591]   <= conv_out_0_591;

    Conv_out[592]   <= conv_out_0_592;

    Conv_out[593]   <= conv_out_0_593;

    Conv_out[594]   <= conv_out_0_594;

    Conv_out[595]   <= conv_out_0_595;

    Conv_out[596]   <= conv_out_0_596;

    Conv_out[597]   <= conv_out_0_597;

    Conv_out[598]   <= conv_out_0_598;

    Conv_out[599]   <= conv_out_0_599;

    Conv_out[600]   <= conv_out_0_600;

    Conv_out[601]   <= conv_out_0_601;

    Conv_out[602]   <= conv_out_0_602;

    Conv_out[603]   <= conv_out_0_603;

    Conv_out[604]   <= conv_out_0_604;

    Conv_out[605]   <= conv_out_0_605;

    Conv_out[606]   <= conv_out_0_606;

    Conv_out[607]   <= conv_out_0_607;

    Conv_out[608]   <= conv_out_0_608;

    Conv_out[609]   <= conv_out_0_609;

    Conv_out[610]   <= conv_out_0_610;

    Conv_out[611]   <= conv_out_0_611;

    Conv_out[612]   <= conv_out_0_612;

    Conv_out[613]   <= conv_out_0_613;

    Conv_out[614]   <= conv_out_0_614;

    Conv_out[615]   <= conv_out_0_615;

    Conv_out[616]   <= conv_out_0_616;

    Conv_out[617]   <= conv_out_0_617;

    Conv_out[618]   <= conv_out_0_618;

    Conv_out[619]   <= conv_out_0_619;

    Conv_out[620]   <= conv_out_0_620;

    Conv_out[621]   <= conv_out_0_621;

    Conv_out[622]   <= conv_out_0_622;

    Conv_out[623]   <= conv_out_0_623;

    Conv_out[624]   <= conv_out_0_624;

    Conv_out[625]   <= conv_out_0_625;

    Conv_out[626]   <= conv_out_0_626;

    Conv_out[627]   <= conv_out_0_627;

    Conv_out[628]   <= conv_out_0_628;

    Conv_out[629]   <= conv_out_0_629;

    Conv_out[630]   <= conv_out_0_630;

    Conv_out[631]   <= conv_out_0_631;

    Conv_out[632]   <= conv_out_0_632;

    Conv_out[633]   <= conv_out_0_633;

    Conv_out[634]   <= conv_out_0_634;

    Conv_out[635]   <= conv_out_0_635;

    Conv_out[636]   <= conv_out_0_636;

    Conv_out[637]   <= conv_out_0_637;

    Conv_out[638]   <= conv_out_0_638;

    Conv_out[639]   <= conv_out_0_639;

    Conv_out[640]   <= conv_out_0_640;

    Conv_out[641]   <= conv_out_0_641;

    Conv_out[642]   <= conv_out_0_642;

    Conv_out[643]   <= conv_out_0_643;

    Conv_out[644]   <= conv_out_0_644;

    Conv_out[645]   <= conv_out_0_645;

    Conv_out[646]   <= conv_out_0_646;

    Conv_out[647]   <= conv_out_0_647;

    Conv_out[648]   <= conv_out_0_648;

    Conv_out[649]   <= conv_out_0_649;

    Conv_out[650]   <= conv_out_0_650;

    Conv_out[651]   <= conv_out_0_651;

    Conv_out[652]   <= conv_out_0_652;

    Conv_out[653]   <= conv_out_0_653;

    Conv_out[654]   <= conv_out_0_654;

    Conv_out[655]   <= conv_out_0_655;

    Conv_out[656]   <= conv_out_0_656;

    Conv_out[657]   <= conv_out_0_657;

    Conv_out[658]   <= conv_out_0_658;

    Conv_out[659]   <= conv_out_0_659;

    Conv_out[660]   <= conv_out_0_660;

    Conv_out[661]   <= conv_out_0_661;

    Conv_out[662]   <= conv_out_0_662;

    Conv_out[663]   <= conv_out_0_663;

    Conv_out[664]   <= conv_out_0_664;

    Conv_out[665]   <= conv_out_0_665;

    Conv_out[666]   <= conv_out_0_666;

    Conv_out[667]   <= conv_out_0_667;

    Conv_out[668]   <= conv_out_0_668;

    Conv_out[669]   <= conv_out_0_669;

    Conv_out[670]   <= conv_out_0_670;

    Conv_out[671]   <= conv_out_0_671;

    Conv_out[672]   <= conv_out_0_672;

    Conv_out[673]   <= conv_out_0_673;

    Conv_out[674]   <= conv_out_0_674;

    Conv_out[675]   <= conv_out_0_675;

    Conv_out[676]   <= conv_out_0_676;

    Conv_out[677]   <= conv_out_0_677;

    Conv_out[678]   <= conv_out_0_678;

    Conv_out[679]   <= conv_out_0_679;

    Conv_out[680]   <= conv_out_0_680;

    Conv_out[681]   <= conv_out_0_681;

    Conv_out[682]   <= conv_out_0_682;

    Conv_out[683]   <= conv_out_0_683;

    Conv_out[684]   <= conv_out_0_684;

    Conv_out[685]   <= conv_out_0_685;

    Conv_out[686]   <= conv_out_0_686;

    Conv_out[687]   <= conv_out_0_687;

    Conv_out[688]   <= conv_out_0_688;

    Conv_out[689]   <= conv_out_0_689;

    Conv_out[690]   <= conv_out_0_690;

    Conv_out[691]   <= conv_out_0_691;

    Conv_out[692]   <= conv_out_0_692;

    Conv_out[693]   <= conv_out_0_693;

    Conv_out[694]   <= conv_out_0_694;

    Conv_out[695]   <= conv_out_0_695;

    Conv_out[696]   <= conv_out_0_696;

    Conv_out[697]   <= conv_out_0_697;

    Conv_out[698]   <= conv_out_0_698;

    Conv_out[699]   <= conv_out_0_699;

    Conv_out[700]   <= conv_out_0_700;

    Conv_out[701]   <= conv_out_0_701;

    Conv_out[702]   <= conv_out_0_702;

    Conv_out[703]   <= conv_out_0_703;

    Conv_out[704]   <= conv_out_0_704;

    Conv_out[705]   <= conv_out_0_705;

    Conv_out[706]   <= conv_out_0_706;

    Conv_out[707]   <= conv_out_0_707;

    Conv_out[708]   <= conv_out_0_708;

    Conv_out[709]   <= conv_out_0_709;

    Conv_out[710]   <= conv_out_0_710;

    Conv_out[711]   <= conv_out_0_711;

    Conv_out[712]   <= conv_out_0_712;

    Conv_out[713]   <= conv_out_0_713;

    Conv_out[714]   <= conv_out_0_714;

    Conv_out[715]   <= conv_out_0_715;

    Conv_out[716]   <= conv_out_0_716;

    Conv_out[717]   <= conv_out_0_717;

    Conv_out[718]   <= conv_out_0_718;

    Conv_out[719]   <= conv_out_0_719;

    Conv_out[720]   <= conv_out_0_720;

    Conv_out[721]   <= conv_out_0_721;

    Conv_out[722]   <= conv_out_0_722;

    Conv_out[723]   <= conv_out_0_723;

    Conv_out[724]   <= conv_out_0_724;

    Conv_out[725]   <= conv_out_0_725;

    Conv_out[726]   <= conv_out_0_726;

    Conv_out[727]   <= conv_out_0_727;

    Conv_out[728]   <= conv_out_0_728;

    Conv_out[729]   <= conv_out_0_729;

    Conv_out[730]   <= conv_out_0_730;

    Conv_out[731]   <= conv_out_0_731;

    Conv_out[732]   <= conv_out_0_732;

    Conv_out[733]   <= conv_out_0_733;

    Conv_out[734]   <= conv_out_0_734;

    Conv_out[735]   <= conv_out_0_735;

    Conv_out[736]   <= conv_out_0_736;

    Conv_out[737]   <= conv_out_0_737;

    Conv_out[738]   <= conv_out_0_738;

    Conv_out[739]   <= conv_out_0_739;

    Conv_out[740]   <= conv_out_0_740;

    Conv_out[741]   <= conv_out_0_741;

    Conv_out[742]   <= conv_out_0_742;

    Conv_out[743]   <= conv_out_0_743;

    Conv_out[744]   <= conv_out_0_744;

    Conv_out[745]   <= conv_out_0_745;

    Conv_out[746]   <= conv_out_0_746;

    Conv_out[747]   <= conv_out_0_747;

    Conv_out[748]   <= conv_out_0_748;

    Conv_out[749]   <= conv_out_0_749;

    Conv_out[750]   <= conv_out_0_750;

    Conv_out[751]   <= conv_out_0_751;

    Conv_out[752]   <= conv_out_0_752;

    Conv_out[753]   <= conv_out_0_753;

    Conv_out[754]   <= conv_out_0_754;

    Conv_out[755]   <= conv_out_0_755;

    Conv_out[756]   <= conv_out_0_756;

    Conv_out[757]   <= conv_out_0_757;

    Conv_out[758]   <= conv_out_0_758;

    Conv_out[759]   <= conv_out_0_759;

    Conv_out[760]   <= conv_out_0_760;

    Conv_out[761]   <= conv_out_0_761;

    Conv_out[762]   <= conv_out_0_762;

    Conv_out[763]   <= conv_out_0_763;

    Conv_out[764]   <= conv_out_0_764;

    Conv_out[765]   <= conv_out_0_765;

    Conv_out[766]   <= conv_out_0_766;

    Conv_out[767]   <= conv_out_0_767;

    Conv_out[768]   <= conv_out_0_768;

    Conv_out[769]   <= conv_out_0_769;

    Conv_out[770]   <= conv_out_0_770;

    Conv_out[771]   <= conv_out_0_771;

    Conv_out[772]   <= conv_out_0_772;

    Conv_out[773]   <= conv_out_0_773;

    Conv_out[774]   <= conv_out_0_774;

    Conv_out[775]   <= conv_out_0_775;

    Conv_out[776]   <= conv_out_0_776;

    Conv_out[777]   <= conv_out_0_777;

    Conv_out[778]   <= conv_out_0_778;

    Conv_out[779]   <= conv_out_0_779;

    Conv_out[780]   <= conv_out_0_780;

    Conv_out[781]   <= conv_out_0_781;

    Conv_out[782]   <= conv_out_0_782;

    Conv_out[783]   <= conv_out_0_783;

    Conv_out[784]   <= conv_out_0_784;

    Conv_out[785]   <= conv_out_0_785;

    Conv_out[786]   <= conv_out_0_786;

    Conv_out[787]   <= conv_out_0_787;

    Conv_out[788]   <= conv_out_0_788;

    Conv_out[789]   <= conv_out_0_789;

    Conv_out[790]   <= conv_out_0_790;

    Conv_out[791]   <= conv_out_0_791;

    Conv_out[792]   <= conv_out_0_792;

    Conv_out[793]   <= conv_out_0_793;

    Conv_out[794]   <= conv_out_0_794;

    Conv_out[795]   <= conv_out_0_795;

    Conv_out[796]   <= conv_out_0_796;

    Conv_out[797]   <= conv_out_0_797;

    Conv_out[798]   <= conv_out_0_798;

    Conv_out[799]   <= conv_out_0_799;

    Conv_out[800]   <= conv_out_0_800;

    Conv_out[801]   <= conv_out_0_801;

    Conv_out[802]   <= conv_out_0_802;

    Conv_out[803]   <= conv_out_0_803;

    Conv_out[804]   <= conv_out_0_804;

    Conv_out[805]   <= conv_out_0_805;

    Conv_out[806]   <= conv_out_0_806;

    Conv_out[807]   <= conv_out_0_807;

    Conv_out[808]   <= conv_out_0_808;

    Conv_out[809]   <= conv_out_0_809;

    Conv_out[810]   <= conv_out_0_810;

    Conv_out[811]   <= conv_out_0_811;

    Conv_out[812]   <= conv_out_0_812;

    Conv_out[813]   <= conv_out_0_813;

    Conv_out[814]   <= conv_out_0_814;

    Conv_out[815]   <= conv_out_0_815;

    Conv_out[816]   <= conv_out_0_816;

    Conv_out[817]   <= conv_out_0_817;

    Conv_out[818]   <= conv_out_0_818;

    Conv_out[819]   <= conv_out_0_819;

    Conv_out[820]   <= conv_out_0_820;

    Conv_out[821]   <= conv_out_0_821;

    Conv_out[822]   <= conv_out_0_822;

    Conv_out[823]   <= conv_out_0_823;

    Conv_out[824]   <= conv_out_0_824;

    Conv_out[825]   <= conv_out_0_825;

    Conv_out[826]   <= conv_out_0_826;

    Conv_out[827]   <= conv_out_0_827;

    Conv_out[828]   <= conv_out_0_828;

    Conv_out[829]   <= conv_out_0_829;

    Conv_out[830]   <= conv_out_0_830;

    Conv_out[831]   <= conv_out_0_831;

    Conv_out[832]   <= conv_out_0_832;

    Conv_out[833]   <= conv_out_0_833;

    Conv_out[834]   <= conv_out_0_834;

    Conv_out[835]   <= conv_out_0_835;

    Conv_out[836]   <= conv_out_0_836;

    Conv_out[837]   <= conv_out_0_837;

    Conv_out[838]   <= conv_out_0_838;

    Conv_out[839]   <= conv_out_0_839;

    Conv_out[840]   <= conv_out_0_840;

    Conv_out[841]   <= conv_out_0_841;

    Conv_out[842]   <= conv_out_0_842;

    Conv_out[843]   <= conv_out_0_843;

    Conv_out[844]   <= conv_out_0_844;

    Conv_out[845]   <= conv_out_0_845;

    Conv_out[846]   <= conv_out_0_846;

    Conv_out[847]   <= conv_out_0_847;

    Conv_out[848]   <= conv_out_0_848;

    Conv_out[849]   <= conv_out_0_849;

    Conv_out[850]   <= conv_out_0_850;

    Conv_out[851]   <= conv_out_0_851;

    Conv_out[852]   <= conv_out_0_852;

    Conv_out[853]   <= conv_out_0_853;

    Conv_out[854]   <= conv_out_0_854;

    Conv_out[855]   <= conv_out_0_855;

    Conv_out[856]   <= conv_out_0_856;

    Conv_out[857]   <= conv_out_0_857;

    Conv_out[858]   <= conv_out_0_858;

    Conv_out[859]   <= conv_out_0_859;

    Conv_out[860]   <= conv_out_0_860;

    Conv_out[861]   <= conv_out_0_861;

    Conv_out[862]   <= conv_out_0_862;

    Conv_out[863]   <= conv_out_0_863;

    Conv_out[864]   <= conv_out_0_864;

    Conv_out[865]   <= conv_out_0_865;

    Conv_out[866]   <= conv_out_0_866;

    Conv_out[867]   <= conv_out_0_867;

    Conv_out[868]   <= conv_out_0_868;

    Conv_out[869]   <= conv_out_0_869;

    Conv_out[870]   <= conv_out_0_870;

    Conv_out[871]   <= conv_out_0_871;

    Conv_out[872]   <= conv_out_0_872;

    Conv_out[873]   <= conv_out_0_873;

    Conv_out[874]   <= conv_out_0_874;

    Conv_out[875]   <= conv_out_0_875;

    Conv_out[876]   <= conv_out_0_876;

    Conv_out[877]   <= conv_out_0_877;

    Conv_out[878]   <= conv_out_0_878;

    Conv_out[879]   <= conv_out_0_879;

    Conv_out[880]   <= conv_out_0_880;

    Conv_out[881]   <= conv_out_0_881;

    Conv_out[882]   <= conv_out_0_882;

    Conv_out[883]   <= conv_out_0_883;

    Conv_out[884]   <= conv_out_0_884;

    Conv_out[885]   <= conv_out_0_885;

    Conv_out[886]   <= conv_out_0_886;

    Conv_out[887]   <= conv_out_0_887;

    Conv_out[888]   <= conv_out_0_888;

    Conv_out[889]   <= conv_out_0_889;

    Conv_out[890]   <= conv_out_0_890;

    Conv_out[891]   <= conv_out_0_891;

    Conv_out[892]   <= conv_out_0_892;

    Conv_out[893]   <= conv_out_0_893;

    Conv_out[894]   <= conv_out_0_894;

    Conv_out[895]   <= conv_out_0_895;

    Conv_out[896]   <= conv_out_0_896;

    Conv_out[897]   <= conv_out_0_897;

    Conv_out[898]   <= conv_out_0_898;

    Conv_out[899]   <= conv_out_0_899;

end

CNN_Single_Layer_2    single0_0(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_0), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_783)
    );

CNN_Single_Layer_2    single0_1(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_1), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_782)
    );

CNN_Single_Layer_2    single0_2(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_2), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_781)
    );

CNN_Single_Layer_2    single0_3(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_3), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_780)
    );

CNN_Single_Layer_2    single0_4(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_4), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_779)
    );

CNN_Single_Layer_2    single0_5(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_5), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_778)
    );

CNN_Single_Layer_2    single0_6(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_6), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_777)
    );

CNN_Single_Layer_2    single0_7(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_7), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_776)
    );

CNN_Single_Layer_2    single0_8(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_8), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_775)
    );

CNN_Single_Layer_2    single0_9(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_9), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_774)
    );

CNN_Single_Layer_2    single0_10(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_10), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_773)
    );

CNN_Single_Layer_2    single0_11(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_11), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_772)
    );

CNN_Single_Layer_2    single0_12(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_12), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_771)
    );

CNN_Single_Layer_2    single0_13(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_13), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_770)
    );

CNN_Single_Layer_2    single0_14(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_14), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_769)
    );

CNN_Single_Layer_2    single0_15(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_15), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_768)
    );

CNN_Single_Layer_2    single0_16(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_16), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_767)
    );

CNN_Single_Layer_2    single0_17(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_17), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_766)
    );

CNN_Single_Layer_2    single0_18(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_18), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_765)
    );

CNN_Single_Layer_2    single0_19(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_19), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_764)
    );

CNN_Single_Layer_2    single0_20(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_20), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_763)
    );

CNN_Single_Layer_2    single0_21(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_21), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_762)
    );

CNN_Single_Layer_2    single0_22(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_22), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_761)
    );

CNN_Single_Layer_2    single0_23(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_23), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_760)
    );

CNN_Single_Layer_2    single0_24(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_24), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_759)
    );

CNN_Single_Layer_2    single0_25(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_25), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_758)
    );

CNN_Single_Layer_2    single0_26(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_26), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_757)
    );

CNN_Single_Layer_2    single0_27(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_27), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_756)
    );

CNN_Single_Layer_2    single0_28(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_28), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_755)
    );

CNN_Single_Layer_2    single0_29(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_29), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_754)
    );

CNN_Single_Layer_2    single0_30(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_30), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_753)
    );

CNN_Single_Layer_2    single0_31(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_31), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_752)
    );

CNN_Single_Layer_2    single0_32(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_32), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_751)
    );

CNN_Single_Layer_2    single0_33(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_33), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_750)
    );

CNN_Single_Layer_2    single0_34(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_34), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_749)
    );

CNN_Single_Layer_2    single0_35(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_35), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_748)
    );

CNN_Single_Layer_2    single0_36(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_36), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_747)
    );

CNN_Single_Layer_2    single0_37(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_37), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_746)
    );

CNN_Single_Layer_2    single0_38(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_38), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_745)
    );

CNN_Single_Layer_2    single0_39(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_39), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_744)
    );

CNN_Single_Layer_2    single0_40(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_40), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_743)
    );

CNN_Single_Layer_2    single0_41(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_41), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_742)
    );

CNN_Single_Layer_2    single0_42(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_42), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_741)
    );

CNN_Single_Layer_2    single0_43(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_43), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_740)
    );

CNN_Single_Layer_2    single0_44(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_44), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_739)
    );

CNN_Single_Layer_2    single0_45(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_45), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_738)
    );

CNN_Single_Layer_2    single0_46(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_46), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_737)
    );

CNN_Single_Layer_2    single0_47(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_47), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_736)
    );

CNN_Single_Layer_2    single0_48(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_48), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_735)
    );

CNN_Single_Layer_2    single0_49(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_49), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_734)
    );

CNN_Single_Layer_2    single0_50(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_50), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_733)
    );

CNN_Single_Layer_2    single0_51(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_51), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_732)
    );

CNN_Single_Layer_2    single0_52(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_52), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_731)
    );

CNN_Single_Layer_2    single0_53(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_53), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_730)
    );

CNN_Single_Layer_2    single0_54(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_54), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_729)
    );

CNN_Single_Layer_2    single0_55(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_55), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_728)
    );

CNN_Single_Layer_2    single0_56(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_56), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_727)
    );

CNN_Single_Layer_2    single0_57(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_57), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_726)
    );

CNN_Single_Layer_2    single0_58(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_58), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_725)
    );

CNN_Single_Layer_2    single0_59(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_59), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_724)
    );

CNN_Single_Layer_2    single0_60(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_60), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_723)
    );

CNN_Single_Layer_2    single0_61(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_61), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_722)
    );

CNN_Single_Layer_2    single0_62(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_62), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_721)
    );

CNN_Single_Layer_2    single0_63(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_63), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_720)
    );

CNN_Single_Layer_2    single0_64(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_64), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_719)
    );

CNN_Single_Layer_2    single0_65(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_65), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_718)
    );

CNN_Single_Layer_2    single0_66(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_66), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_717)
    );

CNN_Single_Layer_2    single0_67(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_67), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_716)
    );

CNN_Single_Layer_2    single0_68(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_68), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_715)
    );

CNN_Single_Layer_2    single0_69(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_69), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_714)
    );

CNN_Single_Layer_2    single0_70(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_70), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_713)
    );

CNN_Single_Layer_2    single0_71(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_71), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_712)
    );

CNN_Single_Layer_2    single0_72(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_72), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_711)
    );

CNN_Single_Layer_2    single0_73(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_73), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_710)
    );

CNN_Single_Layer_2    single0_74(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_74), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_709)
    );

CNN_Single_Layer_2    single0_75(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_75), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_708)
    );

CNN_Single_Layer_2    single0_76(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_76), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_707)
    );

CNN_Single_Layer_2    single0_77(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_77), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_706)
    );

CNN_Single_Layer_2    single0_78(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_78), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_705)
    );

CNN_Single_Layer_2    single0_79(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_79), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_704)
    );

CNN_Single_Layer_2    single0_80(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_80), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_703)
    );

CNN_Single_Layer_2    single0_81(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_81), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_702)
    );

CNN_Single_Layer_2    single0_82(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_82), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_701)
    );

CNN_Single_Layer_2    single0_83(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_83), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_700)
    );

CNN_Single_Layer_2    single0_84(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_84), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_699)
    );

CNN_Single_Layer_2    single0_85(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_85), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_698)
    );

CNN_Single_Layer_2    single0_86(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_86), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_697)
    );

CNN_Single_Layer_2    single0_87(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_87), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_696)
    );

CNN_Single_Layer_2    single0_88(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_88), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_695)
    );

CNN_Single_Layer_2    single0_89(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_89), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_694)
    );

CNN_Single_Layer_2    single0_90(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_90), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_693)
    );

CNN_Single_Layer_2    single0_91(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_91), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_692)
    );

CNN_Single_Layer_2    single0_92(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_92), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_691)
    );

CNN_Single_Layer_2    single0_93(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_93), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_690)
    );

CNN_Single_Layer_2    single0_94(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_94), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_689)
    );

CNN_Single_Layer_2    single0_95(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_95), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_688)
    );

CNN_Single_Layer_2    single0_96(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_96), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_687)
    );

CNN_Single_Layer_2    single0_97(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_97), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_686)
    );

CNN_Single_Layer_2    single0_98(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_98), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_685)
    );

CNN_Single_Layer_2    single0_99(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_99), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_684)
    );

CNN_Single_Layer_2    single0_100(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_100), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_683)
    );

CNN_Single_Layer_2    single0_101(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_101), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_682)
    );

CNN_Single_Layer_2    single0_102(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_102), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_681)
    );

CNN_Single_Layer_2    single0_103(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_103), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_680)
    );

CNN_Single_Layer_2    single0_104(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_104), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_679)
    );

CNN_Single_Layer_2    single0_105(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_105), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_678)
    );

CNN_Single_Layer_2    single0_106(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_106), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_677)
    );

CNN_Single_Layer_2    single0_107(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_107), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_676)
    );

CNN_Single_Layer_2    single0_108(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_108), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_675)
    );

CNN_Single_Layer_2    single0_109(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_109), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_674)
    );

CNN_Single_Layer_2    single0_110(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_110), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_673)
    );

CNN_Single_Layer_2    single0_111(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_111), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_672)
    );

CNN_Single_Layer_2    single0_112(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_112), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_671)
    );

CNN_Single_Layer_2    single0_113(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_113), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_670)
    );

CNN_Single_Layer_2    single0_114(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_114), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_669)
    );

CNN_Single_Layer_2    single0_115(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_115), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_668)
    );

CNN_Single_Layer_2    single0_116(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_116), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_667)
    );

CNN_Single_Layer_2    single0_117(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_117), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_666)
    );

CNN_Single_Layer_2    single0_118(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_118), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_665)
    );

CNN_Single_Layer_2    single0_119(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_119), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_664)
    );

CNN_Single_Layer_2    single0_120(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_120), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_663)
    );

CNN_Single_Layer_2    single0_121(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_121), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_662)
    );

CNN_Single_Layer_2    single0_122(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_122), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_661)
    );

CNN_Single_Layer_2    single0_123(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_123), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_660)
    );

CNN_Single_Layer_2    single0_124(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_124), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_659)
    );

CNN_Single_Layer_2    single0_125(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_125), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_658)
    );

CNN_Single_Layer_2    single0_126(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_126), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_657)
    );

CNN_Single_Layer_2    single0_127(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_127), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_656)
    );

CNN_Single_Layer_2    single0_128(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_128), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_655)
    );

CNN_Single_Layer_2    single0_129(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_129), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_654)
    );

CNN_Single_Layer_2    single0_130(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_130), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_653)
    );

CNN_Single_Layer_2    single0_131(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_131), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_652)
    );

CNN_Single_Layer_2    single0_132(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_132), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_651)
    );

CNN_Single_Layer_2    single0_133(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_133), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_650)
    );

CNN_Single_Layer_2    single0_134(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_134), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_649)
    );

CNN_Single_Layer_2    single0_135(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_135), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_648)
    );

CNN_Single_Layer_2    single0_136(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_136), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_647)
    );

CNN_Single_Layer_2    single0_137(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_137), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_646)
    );

CNN_Single_Layer_2    single0_138(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_138), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_645)
    );

CNN_Single_Layer_2    single0_139(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_139), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_644)
    );

CNN_Single_Layer_2    single0_140(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_140), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_643)
    );

CNN_Single_Layer_2    single0_141(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_141), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_642)
    );

CNN_Single_Layer_2    single0_142(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_142), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_641)
    );

CNN_Single_Layer_2    single0_143(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_143), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_640)
    );

CNN_Single_Layer_2    single0_144(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_144), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_639)
    );

CNN_Single_Layer_2    single0_145(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_145), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_638)
    );

CNN_Single_Layer_2    single0_146(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_146), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_637)
    );

CNN_Single_Layer_2    single0_147(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_147), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_636)
    );

CNN_Single_Layer_2    single0_148(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_148), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_635)
    );

CNN_Single_Layer_2    single0_149(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_149), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_634)
    );

CNN_Single_Layer_2    single0_150(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_150), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_633)
    );

CNN_Single_Layer_2    single0_151(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_151), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_632)
    );

CNN_Single_Layer_2    single0_152(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_152), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_631)
    );

CNN_Single_Layer_2    single0_153(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_153), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_630)
    );

CNN_Single_Layer_2    single0_154(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_154), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_629)
    );

CNN_Single_Layer_2    single0_155(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_155), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_628)
    );

CNN_Single_Layer_2    single0_156(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_156), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_627)
    );

CNN_Single_Layer_2    single0_157(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_157), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_626)
    );

CNN_Single_Layer_2    single0_158(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_158), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_625)
    );

CNN_Single_Layer_2    single0_159(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_159), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_624)
    );

CNN_Single_Layer_2    single0_160(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_160), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_623)
    );

CNN_Single_Layer_2    single0_161(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_161), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_622)
    );

CNN_Single_Layer_2    single0_162(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_162), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_621)
    );

CNN_Single_Layer_2    single0_163(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_163), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_620)
    );

CNN_Single_Layer_2    single0_164(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_164), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_619)
    );

CNN_Single_Layer_2    single0_165(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_165), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_618)
    );

CNN_Single_Layer_2    single0_166(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_166), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_617)
    );

CNN_Single_Layer_2    single0_167(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_167), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_616)
    );

CNN_Single_Layer_2    single0_168(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_168), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_615)
    );

CNN_Single_Layer_2    single0_169(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_169), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_614)
    );

CNN_Single_Layer_2    single0_170(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_170), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_613)
    );

CNN_Single_Layer_2    single0_171(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_171), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_612)
    );

CNN_Single_Layer_2    single0_172(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_172), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_611)
    );

CNN_Single_Layer_2    single0_173(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_173), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_610)
    );

CNN_Single_Layer_2    single0_174(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_174), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_609)
    );

CNN_Single_Layer_2    single0_175(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_175), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_608)
    );

CNN_Single_Layer_2    single0_176(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_176), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_607)
    );

CNN_Single_Layer_2    single0_177(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_177), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_606)
    );

CNN_Single_Layer_2    single0_178(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_178), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_605)
    );

CNN_Single_Layer_2    single0_179(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_179), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_604)
    );

CNN_Single_Layer_2    single0_180(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_180), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_603)
    );

CNN_Single_Layer_2    single0_181(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_181), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_602)
    );

CNN_Single_Layer_2    single0_182(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_182), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_601)
    );

CNN_Single_Layer_2    single0_183(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_183), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_600)
    );

CNN_Single_Layer_2    single0_184(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_184), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_599)
    );

CNN_Single_Layer_2    single0_185(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_185), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_598)
    );

CNN_Single_Layer_2    single0_186(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_186), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_597)
    );

CNN_Single_Layer_2    single0_187(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_187), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_596)
    );

CNN_Single_Layer_2    single0_188(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_188), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_595)
    );

CNN_Single_Layer_2    single0_189(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_189), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_594)
    );

CNN_Single_Layer_2    single0_190(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_190), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_593)
    );

CNN_Single_Layer_2    single0_191(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_191), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_592)
    );

CNN_Single_Layer_2    single0_192(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_192), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_591)
    );

CNN_Single_Layer_2    single0_193(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_193), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_590)
    );

CNN_Single_Layer_2    single0_194(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_194), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_589)
    );

CNN_Single_Layer_2    single0_195(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_195), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_588)
    );

CNN_Single_Layer_2    single0_196(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_196), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_587)
    );

CNN_Single_Layer_2    single0_197(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_197), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_586)
    );

CNN_Single_Layer_2    single0_198(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_198), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_585)
    );

CNN_Single_Layer_2    single0_199(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_199), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_584)
    );

CNN_Single_Layer_2    single0_200(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_200), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_583)
    );

CNN_Single_Layer_2    single0_201(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_201), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_582)
    );

CNN_Single_Layer_2    single0_202(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_202), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_581)
    );

CNN_Single_Layer_2    single0_203(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_203), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_580)
    );

CNN_Single_Layer_2    single0_204(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_204), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_579)
    );

CNN_Single_Layer_2    single0_205(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_205), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_578)
    );

CNN_Single_Layer_2    single0_206(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_206), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_577)
    );

CNN_Single_Layer_2    single0_207(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_207), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_576)
    );

CNN_Single_Layer_2    single0_208(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_208), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_575)
    );

CNN_Single_Layer_2    single0_209(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_209), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_574)
    );

CNN_Single_Layer_2    single0_210(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_210), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_573)
    );

CNN_Single_Layer_2    single0_211(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_211), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_572)
    );

CNN_Single_Layer_2    single0_212(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_212), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_571)
    );

CNN_Single_Layer_2    single0_213(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_213), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_570)
    );

CNN_Single_Layer_2    single0_214(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_214), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_569)
    );

CNN_Single_Layer_2    single0_215(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_215), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_568)
    );

CNN_Single_Layer_2    single0_216(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_216), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_567)
    );

CNN_Single_Layer_2    single0_217(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_217), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_566)
    );

CNN_Single_Layer_2    single0_218(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_218), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_565)
    );

CNN_Single_Layer_2    single0_219(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_219), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_564)
    );

CNN_Single_Layer_2    single0_220(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_220), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_563)
    );

CNN_Single_Layer_2    single0_221(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_221), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_562)
    );

CNN_Single_Layer_2    single0_222(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_222), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_561)
    );

CNN_Single_Layer_2    single0_223(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_223), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_560)
    );

CNN_Single_Layer_2    single0_224(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_224), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_559)
    );

CNN_Single_Layer_2    single0_225(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_225), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_558)
    );

CNN_Single_Layer_2    single0_226(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_226), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_557)
    );

CNN_Single_Layer_2    single0_227(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_227), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_556)
    );

CNN_Single_Layer_2    single0_228(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_228), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_555)
    );

CNN_Single_Layer_2    single0_229(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_229), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_554)
    );

CNN_Single_Layer_2    single0_230(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_230), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_553)
    );

CNN_Single_Layer_2    single0_231(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_231), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_552)
    );

CNN_Single_Layer_2    single0_232(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_232), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_551)
    );

CNN_Single_Layer_2    single0_233(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_233), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_550)
    );

CNN_Single_Layer_2    single0_234(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_234), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_549)
    );

CNN_Single_Layer_2    single0_235(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_235), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_548)
    );

CNN_Single_Layer_2    single0_236(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_236), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_547)
    );

CNN_Single_Layer_2    single0_237(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_237), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_546)
    );

CNN_Single_Layer_2    single0_238(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_238), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_545)
    );

CNN_Single_Layer_2    single0_239(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_239), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_544)
    );

CNN_Single_Layer_2    single0_240(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_240), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_543)
    );

CNN_Single_Layer_2    single0_241(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_241), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_542)
    );

CNN_Single_Layer_2    single0_242(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_242), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_541)
    );

CNN_Single_Layer_2    single0_243(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_243), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_540)
    );

CNN_Single_Layer_2    single0_244(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_244), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_539)
    );

CNN_Single_Layer_2    single0_245(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_245), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_538)
    );

CNN_Single_Layer_2    single0_246(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_246), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_537)
    );

CNN_Single_Layer_2    single0_247(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_247), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_536)
    );

CNN_Single_Layer_2    single0_248(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_248), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_535)
    );

CNN_Single_Layer_2    single0_249(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_249), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_534)
    );

CNN_Single_Layer_2    single0_250(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_250), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_533)
    );

CNN_Single_Layer_2    single0_251(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_251), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_532)
    );

CNN_Single_Layer_2    single0_252(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_252), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_531)
    );

CNN_Single_Layer_2    single0_253(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_253), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_530)
    );

CNN_Single_Layer_2    single0_254(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_254), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_529)
    );

CNN_Single_Layer_2    single0_255(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_255), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_528)
    );

CNN_Single_Layer_2    single0_256(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_256), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_527)
    );

CNN_Single_Layer_2    single0_257(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_257), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_526)
    );

CNN_Single_Layer_2    single0_258(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_258), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_525)
    );

CNN_Single_Layer_2    single0_259(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_259), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_524)
    );

CNN_Single_Layer_2    single0_260(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_260), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_523)
    );

CNN_Single_Layer_2    single0_261(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_261), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_522)
    );

CNN_Single_Layer_2    single0_262(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_262), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_521)
    );

CNN_Single_Layer_2    single0_263(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_263), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_520)
    );

CNN_Single_Layer_2    single0_264(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_264), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_519)
    );

CNN_Single_Layer_2    single0_265(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_265), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_518)
    );

CNN_Single_Layer_2    single0_266(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_266), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_517)
    );

CNN_Single_Layer_2    single0_267(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_267), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_516)
    );

CNN_Single_Layer_2    single0_268(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_268), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_515)
    );

CNN_Single_Layer_2    single0_269(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_269), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_514)
    );

CNN_Single_Layer_2    single0_270(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_270), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_513)
    );

CNN_Single_Layer_2    single0_271(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_271), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_512)
    );

CNN_Single_Layer_2    single0_272(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_272), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_511)
    );

CNN_Single_Layer_2    single0_273(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_273), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_510)
    );

CNN_Single_Layer_2    single0_274(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_274), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_509)
    );

CNN_Single_Layer_2    single0_275(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_275), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_508)
    );

CNN_Single_Layer_2    single0_276(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_276), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_507)
    );

CNN_Single_Layer_2    single0_277(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_277), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_506)
    );

CNN_Single_Layer_2    single0_278(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_278), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_505)
    );

CNN_Single_Layer_2    single0_279(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_279), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_504)
    );

CNN_Single_Layer_2    single0_280(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_280), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_503)
    );

CNN_Single_Layer_2    single0_281(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_281), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_502)
    );

CNN_Single_Layer_2    single0_282(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_282), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_501)
    );

CNN_Single_Layer_2    single0_283(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_283), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_500)
    );

CNN_Single_Layer_2    single0_284(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_284), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_499)
    );

CNN_Single_Layer_2    single0_285(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_285), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_498)
    );

CNN_Single_Layer_2    single0_286(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_286), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_497)
    );

CNN_Single_Layer_2    single0_287(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_287), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_496)
    );

CNN_Single_Layer_2    single0_288(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_288), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_495)
    );

CNN_Single_Layer_2    single0_289(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_289), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_494)
    );

CNN_Single_Layer_2    single0_290(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_290), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_493)
    );

CNN_Single_Layer_2    single0_291(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_291), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_492)
    );

CNN_Single_Layer_2    single0_292(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_292), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_491)
    );

CNN_Single_Layer_2    single0_293(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_293), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_490)
    );

CNN_Single_Layer_2    single0_294(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_294), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_489)
    );

CNN_Single_Layer_2    single0_295(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_295), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_488)
    );

CNN_Single_Layer_2    single0_296(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_296), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_487)
    );

CNN_Single_Layer_2    single0_297(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_297), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_486)
    );

CNN_Single_Layer_2    single0_298(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_298), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_485)
    );

CNN_Single_Layer_2    single0_299(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_299), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_484)
    );

CNN_Single_Layer_2    single0_300(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_300), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_483)
    );

CNN_Single_Layer_2    single0_301(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_301), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_482)
    );

CNN_Single_Layer_2    single0_302(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_302), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_481)
    );

CNN_Single_Layer_2    single0_303(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_303), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_480)
    );

CNN_Single_Layer_2    single0_304(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_304), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_479)
    );

CNN_Single_Layer_2    single0_305(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_305), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_478)
    );

CNN_Single_Layer_2    single0_306(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_306), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_477)
    );

CNN_Single_Layer_2    single0_307(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_307), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_476)
    );

CNN_Single_Layer_2    single0_308(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_308), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_475)
    );

CNN_Single_Layer_2    single0_309(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_309), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_474)
    );

CNN_Single_Layer_2    single0_310(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_310), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_473)
    );

CNN_Single_Layer_2    single0_311(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_311), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_472)
    );

CNN_Single_Layer_2    single0_312(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_312), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_471)
    );

CNN_Single_Layer_2    single0_313(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_313), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_470)
    );

CNN_Single_Layer_2    single0_314(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_314), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_469)
    );

CNN_Single_Layer_2    single0_315(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_315), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_468)
    );

CNN_Single_Layer_2    single0_316(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_316), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_467)
    );

CNN_Single_Layer_2    single0_317(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_317), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_466)
    );

CNN_Single_Layer_2    single0_318(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_318), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_465)
    );

CNN_Single_Layer_2    single0_319(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_319), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_464)
    );

CNN_Single_Layer_2    single0_320(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_320), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_463)
    );

CNN_Single_Layer_2    single0_321(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_321), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_462)
    );

CNN_Single_Layer_2    single0_322(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_322), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_461)
    );

CNN_Single_Layer_2    single0_323(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_323), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_460)
    );

CNN_Single_Layer_2    single0_324(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_324), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_459)
    );

CNN_Single_Layer_2    single0_325(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_325), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_458)
    );

CNN_Single_Layer_2    single0_326(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_326), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_457)
    );

CNN_Single_Layer_2    single0_327(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_327), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_456)
    );

CNN_Single_Layer_2    single0_328(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_328), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_455)
    );

CNN_Single_Layer_2    single0_329(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_329), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_454)
    );

CNN_Single_Layer_2    single0_330(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_330), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_453)
    );

CNN_Single_Layer_2    single0_331(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_331), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_452)
    );

CNN_Single_Layer_2    single0_332(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_332), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_451)
    );

CNN_Single_Layer_2    single0_333(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_333), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_450)
    );

CNN_Single_Layer_2    single0_334(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_334), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_449)
    );

CNN_Single_Layer_2    single0_335(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_335), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_448)
    );

CNN_Single_Layer_2    single0_336(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_336), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_447)
    );

CNN_Single_Layer_2    single0_337(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_337), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_446)
    );

CNN_Single_Layer_2    single0_338(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_338), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_445)
    );

CNN_Single_Layer_2    single0_339(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_339), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_444)
    );

CNN_Single_Layer_2    single0_340(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_340), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_443)
    );

CNN_Single_Layer_2    single0_341(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_341), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_442)
    );

CNN_Single_Layer_2    single0_342(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_342), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_441)
    );

CNN_Single_Layer_2    single0_343(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_343), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_440)
    );

CNN_Single_Layer_2    single0_344(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_344), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_439)
    );

CNN_Single_Layer_2    single0_345(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_345), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_438)
    );

CNN_Single_Layer_2    single0_346(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_346), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_437)
    );

CNN_Single_Layer_2    single0_347(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_347), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_436)
    );

CNN_Single_Layer_2    single0_348(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_348), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_435)
    );

CNN_Single_Layer_2    single0_349(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_349), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_434)
    );

CNN_Single_Layer_2    single0_350(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_350), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_433)
    );

CNN_Single_Layer_2    single0_351(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_351), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_432)
    );

CNN_Single_Layer_2    single0_352(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_352), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_431)
    );

CNN_Single_Layer_2    single0_353(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_353), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_430)
    );

CNN_Single_Layer_2    single0_354(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_354), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_429)
    );

CNN_Single_Layer_2    single0_355(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_355), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_428)
    );

CNN_Single_Layer_2    single0_356(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_356), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_427)
    );

CNN_Single_Layer_2    single0_357(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_357), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_426)
    );

CNN_Single_Layer_2    single0_358(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_358), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_425)
    );

CNN_Single_Layer_2    single0_359(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_359), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_424)
    );

CNN_Single_Layer_2    single0_360(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_360), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_423)
    );

CNN_Single_Layer_2    single0_361(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_361), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_422)
    );

CNN_Single_Layer_2    single0_362(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_362), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_421)
    );

CNN_Single_Layer_2    single0_363(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_363), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_420)
    );

CNN_Single_Layer_2    single0_364(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_364), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_419)
    );

CNN_Single_Layer_2    single0_365(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_365), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_418)
    );

CNN_Single_Layer_2    single0_366(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_366), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_417)
    );

CNN_Single_Layer_2    single0_367(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_367), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_416)
    );

CNN_Single_Layer_2    single0_368(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_368), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_415)
    );

CNN_Single_Layer_2    single0_369(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_369), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_414)
    );

CNN_Single_Layer_2    single0_370(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_370), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_413)
    );

CNN_Single_Layer_2    single0_371(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_371), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_412)
    );

CNN_Single_Layer_2    single0_372(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_372), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_411)
    );

CNN_Single_Layer_2    single0_373(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_373), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_410)
    );

CNN_Single_Layer_2    single0_374(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_374), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_409)
    );

CNN_Single_Layer_2    single0_375(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_375), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_408)
    );

CNN_Single_Layer_2    single0_376(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_376), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_407)
    );

CNN_Single_Layer_2    single0_377(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_377), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_406)
    );

CNN_Single_Layer_2    single0_378(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_378), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_405)
    );

CNN_Single_Layer_2    single0_379(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_379), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_404)
    );

CNN_Single_Layer_2    single0_380(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_380), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_403)
    );

CNN_Single_Layer_2    single0_381(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_381), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_402)
    );

CNN_Single_Layer_2    single0_382(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_382), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_401)
    );

CNN_Single_Layer_2    single0_383(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_383), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_400)
    );

CNN_Single_Layer_2    single0_384(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_384), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_399)
    );

CNN_Single_Layer_2    single0_385(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_385), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_398)
    );

CNN_Single_Layer_2    single0_386(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_386), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_397)
    );

CNN_Single_Layer_2    single0_387(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_387), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_396)
    );

CNN_Single_Layer_2    single0_388(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_388), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_395)
    );

CNN_Single_Layer_2    single0_389(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_389), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_394)
    );

CNN_Single_Layer_2    single0_390(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_390), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_393)
    );

CNN_Single_Layer_2    single0_391(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_391), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_392)
    );

CNN_Single_Layer_2    single0_392(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_392), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_391)
    );

CNN_Single_Layer_2    single0_393(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_393), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_390)
    );

CNN_Single_Layer_2    single0_394(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_394), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_389)
    );

CNN_Single_Layer_2    single0_395(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_395), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_388)
    );

CNN_Single_Layer_2    single0_396(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_396), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_387)
    );

CNN_Single_Layer_2    single0_397(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_397), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_386)
    );

CNN_Single_Layer_2    single0_398(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_398), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_385)
    );

CNN_Single_Layer_2    single0_399(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_399), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_384)
    );

CNN_Single_Layer_2    single0_400(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_400), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_383)
    );

CNN_Single_Layer_2    single0_401(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_401), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_382)
    );

CNN_Single_Layer_2    single0_402(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_402), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_381)
    );

CNN_Single_Layer_2    single0_403(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_403), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_380)
    );

CNN_Single_Layer_2    single0_404(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_404), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_379)
    );

CNN_Single_Layer_2    single0_405(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_405), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_378)
    );

CNN_Single_Layer_2    single0_406(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_406), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_377)
    );

CNN_Single_Layer_2    single0_407(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_407), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_376)
    );

CNN_Single_Layer_2    single0_408(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_408), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_375)
    );

CNN_Single_Layer_2    single0_409(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_409), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_374)
    );

CNN_Single_Layer_2    single0_410(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_410), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_373)
    );

CNN_Single_Layer_2    single0_411(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_411), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_372)
    );

CNN_Single_Layer_2    single0_412(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_412), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_371)
    );

CNN_Single_Layer_2    single0_413(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_413), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_370)
    );

CNN_Single_Layer_2    single0_414(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_414), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_369)
    );

CNN_Single_Layer_2    single0_415(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_415), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_368)
    );

CNN_Single_Layer_2    single0_416(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_416), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_367)
    );

CNN_Single_Layer_2    single0_417(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_417), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_366)
    );

CNN_Single_Layer_2    single0_418(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_418), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_365)
    );

CNN_Single_Layer_2    single0_419(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_419), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_364)
    );

CNN_Single_Layer_2    single0_420(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_420), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_363)
    );

CNN_Single_Layer_2    single0_421(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_421), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_362)
    );

CNN_Single_Layer_2    single0_422(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_422), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_361)
    );

CNN_Single_Layer_2    single0_423(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_423), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_360)
    );

CNN_Single_Layer_2    single0_424(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_424), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_359)
    );

CNN_Single_Layer_2    single0_425(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_425), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_358)
    );

CNN_Single_Layer_2    single0_426(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_426), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_357)
    );

CNN_Single_Layer_2    single0_427(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_427), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_356)
    );

CNN_Single_Layer_2    single0_428(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_428), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_355)
    );

CNN_Single_Layer_2    single0_429(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_429), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_354)
    );

CNN_Single_Layer_2    single0_430(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_430), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_353)
    );

CNN_Single_Layer_2    single0_431(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_431), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_352)
    );

CNN_Single_Layer_2    single0_432(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_432), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_351)
    );

CNN_Single_Layer_2    single0_433(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_433), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_350)
    );

CNN_Single_Layer_2    single0_434(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_434), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_349)
    );

CNN_Single_Layer_2    single0_435(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_435), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_348)
    );

CNN_Single_Layer_2    single0_436(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_436), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_347)
    );

CNN_Single_Layer_2    single0_437(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_437), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_346)
    );

CNN_Single_Layer_2    single0_438(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_438), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_345)
    );

CNN_Single_Layer_2    single0_439(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_439), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_344)
    );

CNN_Single_Layer_2    single0_440(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_440), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_343)
    );

CNN_Single_Layer_2    single0_441(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_441), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_342)
    );

CNN_Single_Layer_2    single0_442(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_442), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_341)
    );

CNN_Single_Layer_2    single0_443(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_443), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_340)
    );

CNN_Single_Layer_2    single0_444(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_444), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_339)
    );

CNN_Single_Layer_2    single0_445(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_445), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_338)
    );

CNN_Single_Layer_2    single0_446(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_446), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_337)
    );

CNN_Single_Layer_2    single0_447(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_447), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_336)
    );

CNN_Single_Layer_2    single0_448(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_448), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_335)
    );

CNN_Single_Layer_2    single0_449(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_449), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_334)
    );

CNN_Single_Layer_2    single0_450(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_450), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_333)
    );

CNN_Single_Layer_2    single0_451(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_451), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_332)
    );

CNN_Single_Layer_2    single0_452(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_452), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_331)
    );

CNN_Single_Layer_2    single0_453(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_453), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_330)
    );

CNN_Single_Layer_2    single0_454(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_454), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_329)
    );

CNN_Single_Layer_2    single0_455(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_455), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_328)
    );

CNN_Single_Layer_2    single0_456(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_456), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_327)
    );

CNN_Single_Layer_2    single0_457(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_457), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_326)
    );

CNN_Single_Layer_2    single0_458(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_458), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_325)
    );

CNN_Single_Layer_2    single0_459(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_459), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_324)
    );

CNN_Single_Layer_2    single0_460(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_460), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_323)
    );

CNN_Single_Layer_2    single0_461(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_461), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_322)
    );

CNN_Single_Layer_2    single0_462(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_462), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_321)
    );

CNN_Single_Layer_2    single0_463(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_463), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_320)
    );

CNN_Single_Layer_2    single0_464(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_464), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_319)
    );

CNN_Single_Layer_2    single0_465(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_465), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_318)
    );

CNN_Single_Layer_2    single0_466(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_466), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_317)
    );

CNN_Single_Layer_2    single0_467(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_467), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_316)
    );

CNN_Single_Layer_2    single0_468(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_468), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_315)
    );

CNN_Single_Layer_2    single0_469(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_469), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_314)
    );

CNN_Single_Layer_2    single0_470(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_470), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_313)
    );

CNN_Single_Layer_2    single0_471(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_471), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_312)
    );

CNN_Single_Layer_2    single0_472(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_472), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_311)
    );

CNN_Single_Layer_2    single0_473(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_473), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_310)
    );

CNN_Single_Layer_2    single0_474(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_474), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_309)
    );

CNN_Single_Layer_2    single0_475(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_475), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_308)
    );

CNN_Single_Layer_2    single0_476(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_476), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_307)
    );

CNN_Single_Layer_2    single0_477(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_477), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_306)
    );

CNN_Single_Layer_2    single0_478(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_478), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_305)
    );

CNN_Single_Layer_2    single0_479(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_479), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_304)
    );

CNN_Single_Layer_2    single0_480(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_480), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_303)
    );

CNN_Single_Layer_2    single0_481(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_481), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_302)
    );

CNN_Single_Layer_2    single0_482(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_482), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_301)
    );

CNN_Single_Layer_2    single0_483(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_483), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_300)
    );

CNN_Single_Layer_2    single0_484(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_484), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_299)
    );

CNN_Single_Layer_2    single0_485(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_485), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_298)
    );

CNN_Single_Layer_2    single0_486(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_486), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_297)
    );

CNN_Single_Layer_2    single0_487(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_487), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_296)
    );

CNN_Single_Layer_2    single0_488(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_488), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_295)
    );

CNN_Single_Layer_2    single0_489(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_489), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_294)
    );

CNN_Single_Layer_2    single0_490(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_490), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_293)
    );

CNN_Single_Layer_2    single0_491(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_491), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_292)
    );

CNN_Single_Layer_2    single0_492(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_492), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_291)
    );

CNN_Single_Layer_2    single0_493(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_493), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_290)
    );

CNN_Single_Layer_2    single0_494(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_494), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_289)
    );

CNN_Single_Layer_2    single0_495(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_495), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_288)
    );

CNN_Single_Layer_2    single0_496(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_496), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_287)
    );

CNN_Single_Layer_2    single0_497(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_497), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_286)
    );

CNN_Single_Layer_2    single0_498(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_498), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_285)
    );

CNN_Single_Layer_2    single0_499(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_499), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_284)
    );

CNN_Single_Layer_2    single0_500(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_500), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_283)
    );

CNN_Single_Layer_2    single0_501(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_501), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_282)
    );

CNN_Single_Layer_2    single0_502(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_502), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_281)
    );

CNN_Single_Layer_2    single0_503(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_503), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_280)
    );

CNN_Single_Layer_2    single0_504(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_504), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_279)
    );

CNN_Single_Layer_2    single0_505(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_505), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_278)
    );

CNN_Single_Layer_2    single0_506(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_506), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_277)
    );

CNN_Single_Layer_2    single0_507(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_507), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_276)
    );

CNN_Single_Layer_2    single0_508(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_508), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_275)
    );

CNN_Single_Layer_2    single0_509(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_509), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_274)
    );

CNN_Single_Layer_2    single0_510(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_510), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_273)
    );

CNN_Single_Layer_2    single0_511(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_511), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_272)
    );

CNN_Single_Layer_2    single0_512(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_512), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_271)
    );

CNN_Single_Layer_2    single0_513(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_513), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_270)
    );

CNN_Single_Layer_2    single0_514(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_514), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_269)
    );

CNN_Single_Layer_2    single0_515(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_515), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_268)
    );

CNN_Single_Layer_2    single0_516(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_516), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_267)
    );

CNN_Single_Layer_2    single0_517(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_517), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_266)
    );

CNN_Single_Layer_2    single0_518(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_518), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_265)
    );

CNN_Single_Layer_2    single0_519(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_519), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_264)
    );

CNN_Single_Layer_2    single0_520(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_520), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_263)
    );

CNN_Single_Layer_2    single0_521(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_521), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_262)
    );

CNN_Single_Layer_2    single0_522(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_522), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_261)
    );

CNN_Single_Layer_2    single0_523(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_523), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_260)
    );

CNN_Single_Layer_2    single0_524(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_524), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_259)
    );

CNN_Single_Layer_2    single0_525(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_525), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_258)
    );

CNN_Single_Layer_2    single0_526(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_526), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_257)
    );

CNN_Single_Layer_2    single0_527(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_527), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_256)
    );

CNN_Single_Layer_2    single0_528(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_528), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_255)
    );

CNN_Single_Layer_2    single0_529(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_529), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_254)
    );

CNN_Single_Layer_2    single0_530(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_530), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_253)
    );

CNN_Single_Layer_2    single0_531(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_531), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_252)
    );

CNN_Single_Layer_2    single0_532(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_532), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_251)
    );

CNN_Single_Layer_2    single0_533(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_533), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_250)
    );

CNN_Single_Layer_2    single0_534(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_534), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_249)
    );

CNN_Single_Layer_2    single0_535(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_535), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_248)
    );

CNN_Single_Layer_2    single0_536(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_536), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_247)
    );

CNN_Single_Layer_2    single0_537(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_537), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_246)
    );

CNN_Single_Layer_2    single0_538(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_538), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_245)
    );

CNN_Single_Layer_2    single0_539(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_539), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_244)
    );

CNN_Single_Layer_2    single0_540(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_540), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_243)
    );

CNN_Single_Layer_2    single0_541(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_541), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_242)
    );

CNN_Single_Layer_2    single0_542(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_542), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_241)
    );

CNN_Single_Layer_2    single0_543(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_543), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_240)
    );

CNN_Single_Layer_2    single0_544(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_544), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_239)
    );

CNN_Single_Layer_2    single0_545(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_545), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_238)
    );

CNN_Single_Layer_2    single0_546(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_546), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_237)
    );

CNN_Single_Layer_2    single0_547(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_547), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_236)
    );

CNN_Single_Layer_2    single0_548(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_548), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_235)
    );

CNN_Single_Layer_2    single0_549(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_549), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_234)
    );

CNN_Single_Layer_2    single0_550(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_550), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_233)
    );

CNN_Single_Layer_2    single0_551(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_551), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_232)
    );

CNN_Single_Layer_2    single0_552(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_552), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_231)
    );

CNN_Single_Layer_2    single0_553(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_553), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_230)
    );

CNN_Single_Layer_2    single0_554(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_554), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_229)
    );

CNN_Single_Layer_2    single0_555(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_555), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_228)
    );

CNN_Single_Layer_2    single0_556(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_556), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_227)
    );

CNN_Single_Layer_2    single0_557(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_557), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_226)
    );

CNN_Single_Layer_2    single0_558(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_558), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_225)
    );

CNN_Single_Layer_2    single0_559(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_559), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_224)
    );

CNN_Single_Layer_2    single0_560(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_560), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_223)
    );

CNN_Single_Layer_2    single0_561(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_561), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_222)
    );

CNN_Single_Layer_2    single0_562(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_562), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_221)
    );

CNN_Single_Layer_2    single0_563(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_563), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_220)
    );

CNN_Single_Layer_2    single0_564(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_564), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_219)
    );

CNN_Single_Layer_2    single0_565(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_565), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_218)
    );

CNN_Single_Layer_2    single0_566(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_566), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_217)
    );

CNN_Single_Layer_2    single0_567(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_567), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_216)
    );

CNN_Single_Layer_2    single0_568(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_568), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_215)
    );

CNN_Single_Layer_2    single0_569(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_569), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_214)
    );

CNN_Single_Layer_2    single0_570(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_570), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_213)
    );

CNN_Single_Layer_2    single0_571(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_571), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_212)
    );

CNN_Single_Layer_2    single0_572(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_572), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_211)
    );

CNN_Single_Layer_2    single0_573(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_573), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_210)
    );

CNN_Single_Layer_2    single0_574(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_574), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_209)
    );

CNN_Single_Layer_2    single0_575(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_575), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_208)
    );

CNN_Single_Layer_2    single0_576(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_576), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_207)
    );

CNN_Single_Layer_2    single0_577(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_577), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_206)
    );

CNN_Single_Layer_2    single0_578(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_578), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_205)
    );

CNN_Single_Layer_2    single0_579(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_579), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_204)
    );

CNN_Single_Layer_2    single0_580(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_580), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_203)
    );

CNN_Single_Layer_2    single0_581(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_581), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_202)
    );

CNN_Single_Layer_2    single0_582(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_582), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_201)
    );

CNN_Single_Layer_2    single0_583(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_583), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_200)
    );

CNN_Single_Layer_2    single0_584(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_584), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_199)
    );

CNN_Single_Layer_2    single0_585(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_585), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_198)
    );

CNN_Single_Layer_2    single0_586(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_586), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_197)
    );

CNN_Single_Layer_2    single0_587(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_587), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_196)
    );

CNN_Single_Layer_2    single0_588(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_588), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_195)
    );

CNN_Single_Layer_2    single0_589(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_589), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_194)
    );

CNN_Single_Layer_2    single0_590(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_590), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_193)
    );

CNN_Single_Layer_2    single0_591(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_591), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_192)
    );

CNN_Single_Layer_2    single0_592(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_592), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_191)
    );

CNN_Single_Layer_2    single0_593(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_593), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_190)
    );

CNN_Single_Layer_2    single0_594(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_594), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_189)
    );

CNN_Single_Layer_2    single0_595(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_595), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_188)
    );

CNN_Single_Layer_2    single0_596(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_596), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_187)
    );

CNN_Single_Layer_2    single0_597(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_597), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_186)
    );

CNN_Single_Layer_2    single0_598(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_598), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_185)
    );

CNN_Single_Layer_2    single0_599(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_599), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_184)
    );

CNN_Single_Layer_2    single0_600(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_600), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_183)
    );

CNN_Single_Layer_2    single0_601(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_601), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_182)
    );

CNN_Single_Layer_2    single0_602(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_602), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_181)
    );

CNN_Single_Layer_2    single0_603(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_603), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_180)
    );

CNN_Single_Layer_2    single0_604(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_604), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_179)
    );

CNN_Single_Layer_2    single0_605(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_605), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_178)
    );

CNN_Single_Layer_2    single0_606(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_606), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_177)
    );

CNN_Single_Layer_2    single0_607(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_607), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_176)
    );

CNN_Single_Layer_2    single0_608(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_608), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_175)
    );

CNN_Single_Layer_2    single0_609(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_609), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_174)
    );

CNN_Single_Layer_2    single0_610(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_610), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_173)
    );

CNN_Single_Layer_2    single0_611(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_611), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_172)
    );

CNN_Single_Layer_2    single0_612(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_612), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_171)
    );

CNN_Single_Layer_2    single0_613(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_613), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_170)
    );

CNN_Single_Layer_2    single0_614(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_614), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_169)
    );

CNN_Single_Layer_2    single0_615(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_615), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_168)
    );

CNN_Single_Layer_2    single0_616(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_616), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_167)
    );

CNN_Single_Layer_2    single0_617(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_617), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_166)
    );

CNN_Single_Layer_2    single0_618(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_618), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_165)
    );

CNN_Single_Layer_2    single0_619(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_619), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_164)
    );

CNN_Single_Layer_2    single0_620(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_620), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_163)
    );

CNN_Single_Layer_2    single0_621(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_621), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_162)
    );

CNN_Single_Layer_2    single0_622(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_622), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_161)
    );

CNN_Single_Layer_2    single0_623(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_623), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_160)
    );

CNN_Single_Layer_2    single0_624(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_624), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_159)
    );

CNN_Single_Layer_2    single0_625(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_625), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_158)
    );

CNN_Single_Layer_2    single0_626(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_626), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_157)
    );

CNN_Single_Layer_2    single0_627(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_627), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_156)
    );

CNN_Single_Layer_2    single0_628(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_628), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_155)
    );

CNN_Single_Layer_2    single0_629(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_629), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_154)
    );

CNN_Single_Layer_2    single0_630(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_630), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_153)
    );

CNN_Single_Layer_2    single0_631(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_631), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_152)
    );

CNN_Single_Layer_2    single0_632(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_632), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_151)
    );

CNN_Single_Layer_2    single0_633(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_633), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_150)
    );

CNN_Single_Layer_2    single0_634(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_634), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_149)
    );

CNN_Single_Layer_2    single0_635(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_635), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_148)
    );

CNN_Single_Layer_2    single0_636(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_636), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_147)
    );

CNN_Single_Layer_2    single0_637(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_637), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_146)
    );

CNN_Single_Layer_2    single0_638(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_638), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_145)
    );

CNN_Single_Layer_2    single0_639(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_639), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_144)
    );

CNN_Single_Layer_2    single0_640(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_640), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_143)
    );

CNN_Single_Layer_2    single0_641(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_641), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_142)
    );

CNN_Single_Layer_2    single0_642(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_642), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_141)
    );

CNN_Single_Layer_2    single0_643(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_643), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_140)
    );

CNN_Single_Layer_2    single0_644(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_644), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_139)
    );

CNN_Single_Layer_2    single0_645(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_645), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_138)
    );

CNN_Single_Layer_2    single0_646(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_646), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_137)
    );

CNN_Single_Layer_2    single0_647(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_647), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_136)
    );

CNN_Single_Layer_2    single0_648(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_648), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_135)
    );

CNN_Single_Layer_2    single0_649(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_649), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_134)
    );

CNN_Single_Layer_2    single0_650(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_650), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_133)
    );

CNN_Single_Layer_2    single0_651(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_651), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_132)
    );

CNN_Single_Layer_2    single0_652(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_652), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_131)
    );

CNN_Single_Layer_2    single0_653(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_653), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_130)
    );

CNN_Single_Layer_2    single0_654(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_654), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_129)
    );

CNN_Single_Layer_2    single0_655(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_655), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_128)
    );

CNN_Single_Layer_2    single0_656(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_656), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_127)
    );

CNN_Single_Layer_2    single0_657(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_657), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_126)
    );

CNN_Single_Layer_2    single0_658(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_658), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_125)
    );

CNN_Single_Layer_2    single0_659(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_659), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_124)
    );

CNN_Single_Layer_2    single0_660(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_660), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_123)
    );

CNN_Single_Layer_2    single0_661(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_661), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_122)
    );

CNN_Single_Layer_2    single0_662(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_662), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_121)
    );

CNN_Single_Layer_2    single0_663(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_663), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_120)
    );

CNN_Single_Layer_2    single0_664(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_664), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_119)
    );

CNN_Single_Layer_2    single0_665(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_665), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_118)
    );

CNN_Single_Layer_2    single0_666(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_666), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_117)
    );

CNN_Single_Layer_2    single0_667(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_667), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_116)
    );

CNN_Single_Layer_2    single0_668(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_668), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_115)
    );

CNN_Single_Layer_2    single0_669(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_669), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_114)
    );

CNN_Single_Layer_2    single0_670(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_670), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_113)
    );

CNN_Single_Layer_2    single0_671(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_671), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_112)
    );

CNN_Single_Layer_2    single0_672(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_672), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_111)
    );

CNN_Single_Layer_2    single0_673(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_673), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_110)
    );

CNN_Single_Layer_2    single0_674(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_674), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_109)
    );

CNN_Single_Layer_2    single0_675(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_675), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_108)
    );

CNN_Single_Layer_2    single0_676(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_676), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_107)
    );

CNN_Single_Layer_2    single0_677(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_677), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_106)
    );

CNN_Single_Layer_2    single0_678(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_678), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_105)
    );

CNN_Single_Layer_2    single0_679(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_679), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_104)
    );

CNN_Single_Layer_2    single0_680(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_680), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_103)
    );

CNN_Single_Layer_2    single0_681(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_681), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_102)
    );

CNN_Single_Layer_2    single0_682(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_682), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_101)
    );

CNN_Single_Layer_2    single0_683(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_683), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_100)
    );

CNN_Single_Layer_2    single0_684(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_684), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_99)
    );

CNN_Single_Layer_2    single0_685(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_685), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_98)
    );

CNN_Single_Layer_2    single0_686(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_686), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_97)
    );

CNN_Single_Layer_2    single0_687(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_687), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_96)
    );

CNN_Single_Layer_2    single0_688(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_688), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_95)
    );

CNN_Single_Layer_2    single0_689(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_689), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_94)
    );

CNN_Single_Layer_2    single0_690(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_690), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_93)
    );

CNN_Single_Layer_2    single0_691(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_691), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_92)
    );

CNN_Single_Layer_2    single0_692(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_692), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_91)
    );

CNN_Single_Layer_2    single0_693(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_693), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_90)
    );

CNN_Single_Layer_2    single0_694(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_694), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_89)
    );

CNN_Single_Layer_2    single0_695(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_695), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_88)
    );

CNN_Single_Layer_2    single0_696(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_696), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_87)
    );

CNN_Single_Layer_2    single0_697(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_697), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_86)
    );

CNN_Single_Layer_2    single0_698(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_698), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_85)
    );

CNN_Single_Layer_2    single0_699(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_699), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_84)
    );

CNN_Single_Layer_2    single0_700(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_700), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_83)
    );

CNN_Single_Layer_2    single0_701(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_701), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_82)
    );

CNN_Single_Layer_2    single0_702(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_702), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_81)
    );

CNN_Single_Layer_2    single0_703(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_703), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_80)
    );

CNN_Single_Layer_2    single0_704(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_704), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_79)
    );

CNN_Single_Layer_2    single0_705(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_705), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_78)
    );

CNN_Single_Layer_2    single0_706(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_706), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_77)
    );

CNN_Single_Layer_2    single0_707(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_707), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_76)
    );

CNN_Single_Layer_2    single0_708(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_708), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_75)
    );

CNN_Single_Layer_2    single0_709(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_709), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_74)
    );

CNN_Single_Layer_2    single0_710(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_710), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_73)
    );

CNN_Single_Layer_2    single0_711(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_711), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_72)
    );

CNN_Single_Layer_2    single0_712(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_712), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_71)
    );

CNN_Single_Layer_2    single0_713(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_713), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_70)
    );

CNN_Single_Layer_2    single0_714(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_714), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_69)
    );

CNN_Single_Layer_2    single0_715(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_715), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_68)
    );

CNN_Single_Layer_2    single0_716(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_716), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_67)
    );

CNN_Single_Layer_2    single0_717(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_717), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_66)
    );

CNN_Single_Layer_2    single0_718(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_718), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_65)
    );

CNN_Single_Layer_2    single0_719(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_719), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_64)
    );

CNN_Single_Layer_2    single0_720(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_720), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_63)
    );

CNN_Single_Layer_2    single0_721(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_721), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_62)
    );

CNN_Single_Layer_2    single0_722(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_722), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_61)
    );

CNN_Single_Layer_2    single0_723(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_723), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_60)
    );

CNN_Single_Layer_2    single0_724(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_724), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_59)
    );

CNN_Single_Layer_2    single0_725(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_725), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_58)
    );

CNN_Single_Layer_2    single0_726(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_726), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_57)
    );

CNN_Single_Layer_2    single0_727(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_727), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_56)
    );

CNN_Single_Layer_2    single0_728(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_728), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_55)
    );

CNN_Single_Layer_2    single0_729(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_729), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_54)
    );

CNN_Single_Layer_2    single0_730(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_730), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_53)
    );

CNN_Single_Layer_2    single0_731(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_731), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_52)
    );

CNN_Single_Layer_2    single0_732(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_732), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_51)
    );

CNN_Single_Layer_2    single0_733(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_733), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_50)
    );

CNN_Single_Layer_2    single0_734(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_734), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_49)
    );

CNN_Single_Layer_2    single0_735(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_735), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_48)
    );

CNN_Single_Layer_2    single0_736(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_736), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_47)
    );

CNN_Single_Layer_2    single0_737(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_737), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_46)
    );

CNN_Single_Layer_2    single0_738(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_738), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_45)
    );

CNN_Single_Layer_2    single0_739(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_739), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_44)
    );

CNN_Single_Layer_2    single0_740(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_740), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_43)
    );

CNN_Single_Layer_2    single0_741(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_741), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_42)
    );

CNN_Single_Layer_2    single0_742(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_742), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_41)
    );

CNN_Single_Layer_2    single0_743(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_743), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_40)
    );

CNN_Single_Layer_2    single0_744(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_744), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_39)
    );

CNN_Single_Layer_2    single0_745(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_745), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_38)
    );

CNN_Single_Layer_2    single0_746(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_746), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_37)
    );

CNN_Single_Layer_2    single0_747(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_747), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_36)
    );

CNN_Single_Layer_2    single0_748(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_748), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_35)
    );

CNN_Single_Layer_2    single0_749(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_749), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_34)
    );

CNN_Single_Layer_2    single0_750(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_750), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_33)
    );

CNN_Single_Layer_2    single0_751(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_751), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_32)
    );

CNN_Single_Layer_2    single0_752(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_752), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_31)
    );

CNN_Single_Layer_2    single0_753(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_753), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_30)
    );

CNN_Single_Layer_2    single0_754(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_754), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_29)
    );

CNN_Single_Layer_2    single0_755(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_755), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_28)
    );

CNN_Single_Layer_2    single0_756(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_756), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_27)
    );

CNN_Single_Layer_2    single0_757(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_757), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_26)
    );

CNN_Single_Layer_2    single0_758(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_758), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_25)
    );

CNN_Single_Layer_2    single0_759(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_759), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_24)
    );

CNN_Single_Layer_2    single0_760(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_760), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_23)
    );

CNN_Single_Layer_2    single0_761(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_761), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_22)
    );

CNN_Single_Layer_2    single0_762(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_762), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_21)
    );

CNN_Single_Layer_2    single0_763(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_763), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_20)
    );

CNN_Single_Layer_2    single0_764(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_764), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_19)
    );

CNN_Single_Layer_2    single0_765(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_765), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_18)
    );

CNN_Single_Layer_2    single0_766(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_766), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_17)
    );

CNN_Single_Layer_2    single0_767(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_767), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_16)
    );

CNN_Single_Layer_2    single0_768(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_768), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_15)
    );

CNN_Single_Layer_2    single0_769(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_769), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_14)
    );

CNN_Single_Layer_2    single0_770(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_770), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_13)
    );

CNN_Single_Layer_2    single0_771(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_771), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_12)
    );

CNN_Single_Layer_2    single0_772(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_772), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_11)
    );

CNN_Single_Layer_2    single0_773(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_773), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_10)
    );

CNN_Single_Layer_2    single0_774(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_774), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_9)
    );

CNN_Single_Layer_2    single0_775(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_775), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_8)
    );

CNN_Single_Layer_2    single0_776(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_776), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_7)
    );

CNN_Single_Layer_2    single0_777(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_777), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_6)
    );

CNN_Single_Layer_2    single0_778(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_778), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_5)
    );

CNN_Single_Layer_2    single0_779(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_779), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_4)
    );

CNN_Single_Layer_2    single0_780(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_780), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_3)
    );

CNN_Single_Layer_2    single0_781(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_781), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_2)
    );

CNN_Single_Layer_2    single0_782(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_782), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_1)
    );

CNN_Single_Layer_2    single0_783(
        .clk(clk), .rst_n(rst_n), .Start(Start), .Image(image_1_783), .Filter(filter), .ReadEn(ReadEn), .ConvResult(conv_out_1_0)
    );



    always @(*) begin
    Conv_out_2[0]   <= conv_out_1_0;

    Conv_out_2[1]   <= conv_out_1_1;

    Conv_out_2[2]   <= conv_out_1_2;

    Conv_out_2[3]   <= conv_out_1_3;

    Conv_out_2[4]   <= conv_out_1_4;

    Conv_out_2[5]   <= conv_out_1_5;

    Conv_out_2[6]   <= conv_out_1_6;

    Conv_out_2[7]   <= conv_out_1_7;

    Conv_out_2[8]   <= conv_out_1_8;

    Conv_out_2[9]   <= conv_out_1_9;

    Conv_out_2[10]   <= conv_out_1_10;

    Conv_out_2[11]   <= conv_out_1_11;

    Conv_out_2[12]   <= conv_out_1_12;

    Conv_out_2[13]   <= conv_out_1_13;

    Conv_out_2[14]   <= conv_out_1_14;

    Conv_out_2[15]   <= conv_out_1_15;

    Conv_out_2[16]   <= conv_out_1_16;

    Conv_out_2[17]   <= conv_out_1_17;

    Conv_out_2[18]   <= conv_out_1_18;

    Conv_out_2[19]   <= conv_out_1_19;

    Conv_out_2[20]   <= conv_out_1_20;

    Conv_out_2[21]   <= conv_out_1_21;

    Conv_out_2[22]   <= conv_out_1_22;

    Conv_out_2[23]   <= conv_out_1_23;

    Conv_out_2[24]   <= conv_out_1_24;

    Conv_out_2[25]   <= conv_out_1_25;

    Conv_out_2[26]   <= conv_out_1_26;

    Conv_out_2[27]   <= conv_out_1_27;

    Conv_out_2[28]   <= conv_out_1_28;

    Conv_out_2[29]   <= conv_out_1_29;

    Conv_out_2[30]   <= conv_out_1_30;

    Conv_out_2[31]   <= conv_out_1_31;

    Conv_out_2[32]   <= conv_out_1_32;

    Conv_out_2[33]   <= conv_out_1_33;

    Conv_out_2[34]   <= conv_out_1_34;

    Conv_out_2[35]   <= conv_out_1_35;

    Conv_out_2[36]   <= conv_out_1_36;

    Conv_out_2[37]   <= conv_out_1_37;

    Conv_out_2[38]   <= conv_out_1_38;

    Conv_out_2[39]   <= conv_out_1_39;

    Conv_out_2[40]   <= conv_out_1_40;

    Conv_out_2[41]   <= conv_out_1_41;

    Conv_out_2[42]   <= conv_out_1_42;

    Conv_out_2[43]   <= conv_out_1_43;

    Conv_out_2[44]   <= conv_out_1_44;

    Conv_out_2[45]   <= conv_out_1_45;

    Conv_out_2[46]   <= conv_out_1_46;

    Conv_out_2[47]   <= conv_out_1_47;

    Conv_out_2[48]   <= conv_out_1_48;

    Conv_out_2[49]   <= conv_out_1_49;

    Conv_out_2[50]   <= conv_out_1_50;

    Conv_out_2[51]   <= conv_out_1_51;

    Conv_out_2[52]   <= conv_out_1_52;

    Conv_out_2[53]   <= conv_out_1_53;

    Conv_out_2[54]   <= conv_out_1_54;

    Conv_out_2[55]   <= conv_out_1_55;

    Conv_out_2[56]   <= conv_out_1_56;

    Conv_out_2[57]   <= conv_out_1_57;

    Conv_out_2[58]   <= conv_out_1_58;

    Conv_out_2[59]   <= conv_out_1_59;

    Conv_out_2[60]   <= conv_out_1_60;

    Conv_out_2[61]   <= conv_out_1_61;

    Conv_out_2[62]   <= conv_out_1_62;

    Conv_out_2[63]   <= conv_out_1_63;

    Conv_out_2[64]   <= conv_out_1_64;

    Conv_out_2[65]   <= conv_out_1_65;

    Conv_out_2[66]   <= conv_out_1_66;

    Conv_out_2[67]   <= conv_out_1_67;

    Conv_out_2[68]   <= conv_out_1_68;

    Conv_out_2[69]   <= conv_out_1_69;

    Conv_out_2[70]   <= conv_out_1_70;

    Conv_out_2[71]   <= conv_out_1_71;

    Conv_out_2[72]   <= conv_out_1_72;

    Conv_out_2[73]   <= conv_out_1_73;

    Conv_out_2[74]   <= conv_out_1_74;

    Conv_out_2[75]   <= conv_out_1_75;

    Conv_out_2[76]   <= conv_out_1_76;

    Conv_out_2[77]   <= conv_out_1_77;

    Conv_out_2[78]   <= conv_out_1_78;

    Conv_out_2[79]   <= conv_out_1_79;

    Conv_out_2[80]   <= conv_out_1_80;

    Conv_out_2[81]   <= conv_out_1_81;

    Conv_out_2[82]   <= conv_out_1_82;

    Conv_out_2[83]   <= conv_out_1_83;

    Conv_out_2[84]   <= conv_out_1_84;

    Conv_out_2[85]   <= conv_out_1_85;

    Conv_out_2[86]   <= conv_out_1_86;

    Conv_out_2[87]   <= conv_out_1_87;

    Conv_out_2[88]   <= conv_out_1_88;

    Conv_out_2[89]   <= conv_out_1_89;

    Conv_out_2[90]   <= conv_out_1_90;

    Conv_out_2[91]   <= conv_out_1_91;

    Conv_out_2[92]   <= conv_out_1_92;

    Conv_out_2[93]   <= conv_out_1_93;

    Conv_out_2[94]   <= conv_out_1_94;

    Conv_out_2[95]   <= conv_out_1_95;

    Conv_out_2[96]   <= conv_out_1_96;

    Conv_out_2[97]   <= conv_out_1_97;

    Conv_out_2[98]   <= conv_out_1_98;

    Conv_out_2[99]   <= conv_out_1_99;

    Conv_out_2[100]   <= conv_out_1_100;

    Conv_out_2[101]   <= conv_out_1_101;

    Conv_out_2[102]   <= conv_out_1_102;

    Conv_out_2[103]   <= conv_out_1_103;

    Conv_out_2[104]   <= conv_out_1_104;

    Conv_out_2[105]   <= conv_out_1_105;

    Conv_out_2[106]   <= conv_out_1_106;

    Conv_out_2[107]   <= conv_out_1_107;

    Conv_out_2[108]   <= conv_out_1_108;

    Conv_out_2[109]   <= conv_out_1_109;

    Conv_out_2[110]   <= conv_out_1_110;

    Conv_out_2[111]   <= conv_out_1_111;

    Conv_out_2[112]   <= conv_out_1_112;

    Conv_out_2[113]   <= conv_out_1_113;

    Conv_out_2[114]   <= conv_out_1_114;

    Conv_out_2[115]   <= conv_out_1_115;

    Conv_out_2[116]   <= conv_out_1_116;

    Conv_out_2[117]   <= conv_out_1_117;

    Conv_out_2[118]   <= conv_out_1_118;

    Conv_out_2[119]   <= conv_out_1_119;

    Conv_out_2[120]   <= conv_out_1_120;

    Conv_out_2[121]   <= conv_out_1_121;

    Conv_out_2[122]   <= conv_out_1_122;

    Conv_out_2[123]   <= conv_out_1_123;

    Conv_out_2[124]   <= conv_out_1_124;

    Conv_out_2[125]   <= conv_out_1_125;

    Conv_out_2[126]   <= conv_out_1_126;

    Conv_out_2[127]   <= conv_out_1_127;

    Conv_out_2[128]   <= conv_out_1_128;

    Conv_out_2[129]   <= conv_out_1_129;

    Conv_out_2[130]   <= conv_out_1_130;

    Conv_out_2[131]   <= conv_out_1_131;

    Conv_out_2[132]   <= conv_out_1_132;

    Conv_out_2[133]   <= conv_out_1_133;

    Conv_out_2[134]   <= conv_out_1_134;

    Conv_out_2[135]   <= conv_out_1_135;

    Conv_out_2[136]   <= conv_out_1_136;

    Conv_out_2[137]   <= conv_out_1_137;

    Conv_out_2[138]   <= conv_out_1_138;

    Conv_out_2[139]   <= conv_out_1_139;

    Conv_out_2[140]   <= conv_out_1_140;

    Conv_out_2[141]   <= conv_out_1_141;

    Conv_out_2[142]   <= conv_out_1_142;

    Conv_out_2[143]   <= conv_out_1_143;

    Conv_out_2[144]   <= conv_out_1_144;

    Conv_out_2[145]   <= conv_out_1_145;

    Conv_out_2[146]   <= conv_out_1_146;

    Conv_out_2[147]   <= conv_out_1_147;

    Conv_out_2[148]   <= conv_out_1_148;

    Conv_out_2[149]   <= conv_out_1_149;

    Conv_out_2[150]   <= conv_out_1_150;

    Conv_out_2[151]   <= conv_out_1_151;

    Conv_out_2[152]   <= conv_out_1_152;

    Conv_out_2[153]   <= conv_out_1_153;

    Conv_out_2[154]   <= conv_out_1_154;

    Conv_out_2[155]   <= conv_out_1_155;

    Conv_out_2[156]   <= conv_out_1_156;

    Conv_out_2[157]   <= conv_out_1_157;

    Conv_out_2[158]   <= conv_out_1_158;

    Conv_out_2[159]   <= conv_out_1_159;

    Conv_out_2[160]   <= conv_out_1_160;

    Conv_out_2[161]   <= conv_out_1_161;

    Conv_out_2[162]   <= conv_out_1_162;

    Conv_out_2[163]   <= conv_out_1_163;

    Conv_out_2[164]   <= conv_out_1_164;

    Conv_out_2[165]   <= conv_out_1_165;

    Conv_out_2[166]   <= conv_out_1_166;

    Conv_out_2[167]   <= conv_out_1_167;

    Conv_out_2[168]   <= conv_out_1_168;

    Conv_out_2[169]   <= conv_out_1_169;

    Conv_out_2[170]   <= conv_out_1_170;

    Conv_out_2[171]   <= conv_out_1_171;

    Conv_out_2[172]   <= conv_out_1_172;

    Conv_out_2[173]   <= conv_out_1_173;

    Conv_out_2[174]   <= conv_out_1_174;

    Conv_out_2[175]   <= conv_out_1_175;

    Conv_out_2[176]   <= conv_out_1_176;

    Conv_out_2[177]   <= conv_out_1_177;

    Conv_out_2[178]   <= conv_out_1_178;

    Conv_out_2[179]   <= conv_out_1_179;

    Conv_out_2[180]   <= conv_out_1_180;

    Conv_out_2[181]   <= conv_out_1_181;

    Conv_out_2[182]   <= conv_out_1_182;

    Conv_out_2[183]   <= conv_out_1_183;

    Conv_out_2[184]   <= conv_out_1_184;

    Conv_out_2[185]   <= conv_out_1_185;

    Conv_out_2[186]   <= conv_out_1_186;

    Conv_out_2[187]   <= conv_out_1_187;

    Conv_out_2[188]   <= conv_out_1_188;

    Conv_out_2[189]   <= conv_out_1_189;

    Conv_out_2[190]   <= conv_out_1_190;

    Conv_out_2[191]   <= conv_out_1_191;

    Conv_out_2[192]   <= conv_out_1_192;

    Conv_out_2[193]   <= conv_out_1_193;

    Conv_out_2[194]   <= conv_out_1_194;

    Conv_out_2[195]   <= conv_out_1_195;

    Conv_out_2[196]   <= conv_out_1_196;

    Conv_out_2[197]   <= conv_out_1_197;

    Conv_out_2[198]   <= conv_out_1_198;

    Conv_out_2[199]   <= conv_out_1_199;

    Conv_out_2[200]   <= conv_out_1_200;

    Conv_out_2[201]   <= conv_out_1_201;

    Conv_out_2[202]   <= conv_out_1_202;

    Conv_out_2[203]   <= conv_out_1_203;

    Conv_out_2[204]   <= conv_out_1_204;

    Conv_out_2[205]   <= conv_out_1_205;

    Conv_out_2[206]   <= conv_out_1_206;

    Conv_out_2[207]   <= conv_out_1_207;

    Conv_out_2[208]   <= conv_out_1_208;

    Conv_out_2[209]   <= conv_out_1_209;

    Conv_out_2[210]   <= conv_out_1_210;

    Conv_out_2[211]   <= conv_out_1_211;

    Conv_out_2[212]   <= conv_out_1_212;

    Conv_out_2[213]   <= conv_out_1_213;

    Conv_out_2[214]   <= conv_out_1_214;

    Conv_out_2[215]   <= conv_out_1_215;

    Conv_out_2[216]   <= conv_out_1_216;

    Conv_out_2[217]   <= conv_out_1_217;

    Conv_out_2[218]   <= conv_out_1_218;

    Conv_out_2[219]   <= conv_out_1_219;

    Conv_out_2[220]   <= conv_out_1_220;

    Conv_out_2[221]   <= conv_out_1_221;

    Conv_out_2[222]   <= conv_out_1_222;

    Conv_out_2[223]   <= conv_out_1_223;

    Conv_out_2[224]   <= conv_out_1_224;

    Conv_out_2[225]   <= conv_out_1_225;

    Conv_out_2[226]   <= conv_out_1_226;

    Conv_out_2[227]   <= conv_out_1_227;

    Conv_out_2[228]   <= conv_out_1_228;

    Conv_out_2[229]   <= conv_out_1_229;

    Conv_out_2[230]   <= conv_out_1_230;

    Conv_out_2[231]   <= conv_out_1_231;

    Conv_out_2[232]   <= conv_out_1_232;

    Conv_out_2[233]   <= conv_out_1_233;

    Conv_out_2[234]   <= conv_out_1_234;

    Conv_out_2[235]   <= conv_out_1_235;

    Conv_out_2[236]   <= conv_out_1_236;

    Conv_out_2[237]   <= conv_out_1_237;

    Conv_out_2[238]   <= conv_out_1_238;

    Conv_out_2[239]   <= conv_out_1_239;

    Conv_out_2[240]   <= conv_out_1_240;

    Conv_out_2[241]   <= conv_out_1_241;

    Conv_out_2[242]   <= conv_out_1_242;

    Conv_out_2[243]   <= conv_out_1_243;

    Conv_out_2[244]   <= conv_out_1_244;

    Conv_out_2[245]   <= conv_out_1_245;

    Conv_out_2[246]   <= conv_out_1_246;

    Conv_out_2[247]   <= conv_out_1_247;

    Conv_out_2[248]   <= conv_out_1_248;

    Conv_out_2[249]   <= conv_out_1_249;

    Conv_out_2[250]   <= conv_out_1_250;

    Conv_out_2[251]   <= conv_out_1_251;

    Conv_out_2[252]   <= conv_out_1_252;

    Conv_out_2[253]   <= conv_out_1_253;

    Conv_out_2[254]   <= conv_out_1_254;

    Conv_out_2[255]   <= conv_out_1_255;

    Conv_out_2[256]   <= conv_out_1_256;

    Conv_out_2[257]   <= conv_out_1_257;

    Conv_out_2[258]   <= conv_out_1_258;

    Conv_out_2[259]   <= conv_out_1_259;

    Conv_out_2[260]   <= conv_out_1_260;

    Conv_out_2[261]   <= conv_out_1_261;

    Conv_out_2[262]   <= conv_out_1_262;

    Conv_out_2[263]   <= conv_out_1_263;

    Conv_out_2[264]   <= conv_out_1_264;

    Conv_out_2[265]   <= conv_out_1_265;

    Conv_out_2[266]   <= conv_out_1_266;

    Conv_out_2[267]   <= conv_out_1_267;

    Conv_out_2[268]   <= conv_out_1_268;

    Conv_out_2[269]   <= conv_out_1_269;

    Conv_out_2[270]   <= conv_out_1_270;

    Conv_out_2[271]   <= conv_out_1_271;

    Conv_out_2[272]   <= conv_out_1_272;

    Conv_out_2[273]   <= conv_out_1_273;

    Conv_out_2[274]   <= conv_out_1_274;

    Conv_out_2[275]   <= conv_out_1_275;

    Conv_out_2[276]   <= conv_out_1_276;

    Conv_out_2[277]   <= conv_out_1_277;

    Conv_out_2[278]   <= conv_out_1_278;

    Conv_out_2[279]   <= conv_out_1_279;

    Conv_out_2[280]   <= conv_out_1_280;

    Conv_out_2[281]   <= conv_out_1_281;

    Conv_out_2[282]   <= conv_out_1_282;

    Conv_out_2[283]   <= conv_out_1_283;

    Conv_out_2[284]   <= conv_out_1_284;

    Conv_out_2[285]   <= conv_out_1_285;

    Conv_out_2[286]   <= conv_out_1_286;

    Conv_out_2[287]   <= conv_out_1_287;

    Conv_out_2[288]   <= conv_out_1_288;

    Conv_out_2[289]   <= conv_out_1_289;

    Conv_out_2[290]   <= conv_out_1_290;

    Conv_out_2[291]   <= conv_out_1_291;

    Conv_out_2[292]   <= conv_out_1_292;

    Conv_out_2[293]   <= conv_out_1_293;

    Conv_out_2[294]   <= conv_out_1_294;

    Conv_out_2[295]   <= conv_out_1_295;

    Conv_out_2[296]   <= conv_out_1_296;

    Conv_out_2[297]   <= conv_out_1_297;

    Conv_out_2[298]   <= conv_out_1_298;

    Conv_out_2[299]   <= conv_out_1_299;

    Conv_out_2[300]   <= conv_out_1_300;

    Conv_out_2[301]   <= conv_out_1_301;

    Conv_out_2[302]   <= conv_out_1_302;

    Conv_out_2[303]   <= conv_out_1_303;

    Conv_out_2[304]   <= conv_out_1_304;

    Conv_out_2[305]   <= conv_out_1_305;

    Conv_out_2[306]   <= conv_out_1_306;

    Conv_out_2[307]   <= conv_out_1_307;

    Conv_out_2[308]   <= conv_out_1_308;

    Conv_out_2[309]   <= conv_out_1_309;

    Conv_out_2[310]   <= conv_out_1_310;

    Conv_out_2[311]   <= conv_out_1_311;

    Conv_out_2[312]   <= conv_out_1_312;

    Conv_out_2[313]   <= conv_out_1_313;

    Conv_out_2[314]   <= conv_out_1_314;

    Conv_out_2[315]   <= conv_out_1_315;

    Conv_out_2[316]   <= conv_out_1_316;

    Conv_out_2[317]   <= conv_out_1_317;

    Conv_out_2[318]   <= conv_out_1_318;

    Conv_out_2[319]   <= conv_out_1_319;

    Conv_out_2[320]   <= conv_out_1_320;

    Conv_out_2[321]   <= conv_out_1_321;

    Conv_out_2[322]   <= conv_out_1_322;

    Conv_out_2[323]   <= conv_out_1_323;

    Conv_out_2[324]   <= conv_out_1_324;

    Conv_out_2[325]   <= conv_out_1_325;

    Conv_out_2[326]   <= conv_out_1_326;

    Conv_out_2[327]   <= conv_out_1_327;

    Conv_out_2[328]   <= conv_out_1_328;

    Conv_out_2[329]   <= conv_out_1_329;

    Conv_out_2[330]   <= conv_out_1_330;

    Conv_out_2[331]   <= conv_out_1_331;

    Conv_out_2[332]   <= conv_out_1_332;

    Conv_out_2[333]   <= conv_out_1_333;

    Conv_out_2[334]   <= conv_out_1_334;

    Conv_out_2[335]   <= conv_out_1_335;

    Conv_out_2[336]   <= conv_out_1_336;

    Conv_out_2[337]   <= conv_out_1_337;

    Conv_out_2[338]   <= conv_out_1_338;

    Conv_out_2[339]   <= conv_out_1_339;

    Conv_out_2[340]   <= conv_out_1_340;

    Conv_out_2[341]   <= conv_out_1_341;

    Conv_out_2[342]   <= conv_out_1_342;

    Conv_out_2[343]   <= conv_out_1_343;

    Conv_out_2[344]   <= conv_out_1_344;

    Conv_out_2[345]   <= conv_out_1_345;

    Conv_out_2[346]   <= conv_out_1_346;

    Conv_out_2[347]   <= conv_out_1_347;

    Conv_out_2[348]   <= conv_out_1_348;

    Conv_out_2[349]   <= conv_out_1_349;

    Conv_out_2[350]   <= conv_out_1_350;

    Conv_out_2[351]   <= conv_out_1_351;

    Conv_out_2[352]   <= conv_out_1_352;

    Conv_out_2[353]   <= conv_out_1_353;

    Conv_out_2[354]   <= conv_out_1_354;

    Conv_out_2[355]   <= conv_out_1_355;

    Conv_out_2[356]   <= conv_out_1_356;

    Conv_out_2[357]   <= conv_out_1_357;

    Conv_out_2[358]   <= conv_out_1_358;

    Conv_out_2[359]   <= conv_out_1_359;

    Conv_out_2[360]   <= conv_out_1_360;

    Conv_out_2[361]   <= conv_out_1_361;

    Conv_out_2[362]   <= conv_out_1_362;

    Conv_out_2[363]   <= conv_out_1_363;

    Conv_out_2[364]   <= conv_out_1_364;

    Conv_out_2[365]   <= conv_out_1_365;

    Conv_out_2[366]   <= conv_out_1_366;

    Conv_out_2[367]   <= conv_out_1_367;

    Conv_out_2[368]   <= conv_out_1_368;

    Conv_out_2[369]   <= conv_out_1_369;

    Conv_out_2[370]   <= conv_out_1_370;

    Conv_out_2[371]   <= conv_out_1_371;

    Conv_out_2[372]   <= conv_out_1_372;

    Conv_out_2[373]   <= conv_out_1_373;

    Conv_out_2[374]   <= conv_out_1_374;

    Conv_out_2[375]   <= conv_out_1_375;

    Conv_out_2[376]   <= conv_out_1_376;

    Conv_out_2[377]   <= conv_out_1_377;

    Conv_out_2[378]   <= conv_out_1_378;

    Conv_out_2[379]   <= conv_out_1_379;

    Conv_out_2[380]   <= conv_out_1_380;

    Conv_out_2[381]   <= conv_out_1_381;

    Conv_out_2[382]   <= conv_out_1_382;

    Conv_out_2[383]   <= conv_out_1_383;

    Conv_out_2[384]   <= conv_out_1_384;

    Conv_out_2[385]   <= conv_out_1_385;

    Conv_out_2[386]   <= conv_out_1_386;

    Conv_out_2[387]   <= conv_out_1_387;

    Conv_out_2[388]   <= conv_out_1_388;

    Conv_out_2[389]   <= conv_out_1_389;

    Conv_out_2[390]   <= conv_out_1_390;

    Conv_out_2[391]   <= conv_out_1_391;

    Conv_out_2[392]   <= conv_out_1_392;

    Conv_out_2[393]   <= conv_out_1_393;

    Conv_out_2[394]   <= conv_out_1_394;

    Conv_out_2[395]   <= conv_out_1_395;

    Conv_out_2[396]   <= conv_out_1_396;

    Conv_out_2[397]   <= conv_out_1_397;

    Conv_out_2[398]   <= conv_out_1_398;

    Conv_out_2[399]   <= conv_out_1_399;

    Conv_out_2[400]   <= conv_out_1_400;

    Conv_out_2[401]   <= conv_out_1_401;

    Conv_out_2[402]   <= conv_out_1_402;

    Conv_out_2[403]   <= conv_out_1_403;

    Conv_out_2[404]   <= conv_out_1_404;

    Conv_out_2[405]   <= conv_out_1_405;

    Conv_out_2[406]   <= conv_out_1_406;

    Conv_out_2[407]   <= conv_out_1_407;

    Conv_out_2[408]   <= conv_out_1_408;

    Conv_out_2[409]   <= conv_out_1_409;

    Conv_out_2[410]   <= conv_out_1_410;

    Conv_out_2[411]   <= conv_out_1_411;

    Conv_out_2[412]   <= conv_out_1_412;

    Conv_out_2[413]   <= conv_out_1_413;

    Conv_out_2[414]   <= conv_out_1_414;

    Conv_out_2[415]   <= conv_out_1_415;

    Conv_out_2[416]   <= conv_out_1_416;

    Conv_out_2[417]   <= conv_out_1_417;

    Conv_out_2[418]   <= conv_out_1_418;

    Conv_out_2[419]   <= conv_out_1_419;

    Conv_out_2[420]   <= conv_out_1_420;

    Conv_out_2[421]   <= conv_out_1_421;

    Conv_out_2[422]   <= conv_out_1_422;

    Conv_out_2[423]   <= conv_out_1_423;

    Conv_out_2[424]   <= conv_out_1_424;

    Conv_out_2[425]   <= conv_out_1_425;

    Conv_out_2[426]   <= conv_out_1_426;

    Conv_out_2[427]   <= conv_out_1_427;

    Conv_out_2[428]   <= conv_out_1_428;

    Conv_out_2[429]   <= conv_out_1_429;

    Conv_out_2[430]   <= conv_out_1_430;

    Conv_out_2[431]   <= conv_out_1_431;

    Conv_out_2[432]   <= conv_out_1_432;

    Conv_out_2[433]   <= conv_out_1_433;

    Conv_out_2[434]   <= conv_out_1_434;

    Conv_out_2[435]   <= conv_out_1_435;

    Conv_out_2[436]   <= conv_out_1_436;

    Conv_out_2[437]   <= conv_out_1_437;

    Conv_out_2[438]   <= conv_out_1_438;

    Conv_out_2[439]   <= conv_out_1_439;

    Conv_out_2[440]   <= conv_out_1_440;

    Conv_out_2[441]   <= conv_out_1_441;

    Conv_out_2[442]   <= conv_out_1_442;

    Conv_out_2[443]   <= conv_out_1_443;

    Conv_out_2[444]   <= conv_out_1_444;

    Conv_out_2[445]   <= conv_out_1_445;

    Conv_out_2[446]   <= conv_out_1_446;

    Conv_out_2[447]   <= conv_out_1_447;

    Conv_out_2[448]   <= conv_out_1_448;

    Conv_out_2[449]   <= conv_out_1_449;

    Conv_out_2[450]   <= conv_out_1_450;

    Conv_out_2[451]   <= conv_out_1_451;

    Conv_out_2[452]   <= conv_out_1_452;

    Conv_out_2[453]   <= conv_out_1_453;

    Conv_out_2[454]   <= conv_out_1_454;

    Conv_out_2[455]   <= conv_out_1_455;

    Conv_out_2[456]   <= conv_out_1_456;

    Conv_out_2[457]   <= conv_out_1_457;

    Conv_out_2[458]   <= conv_out_1_458;

    Conv_out_2[459]   <= conv_out_1_459;

    Conv_out_2[460]   <= conv_out_1_460;

    Conv_out_2[461]   <= conv_out_1_461;

    Conv_out_2[462]   <= conv_out_1_462;

    Conv_out_2[463]   <= conv_out_1_463;

    Conv_out_2[464]   <= conv_out_1_464;

    Conv_out_2[465]   <= conv_out_1_465;

    Conv_out_2[466]   <= conv_out_1_466;

    Conv_out_2[467]   <= conv_out_1_467;

    Conv_out_2[468]   <= conv_out_1_468;

    Conv_out_2[469]   <= conv_out_1_469;

    Conv_out_2[470]   <= conv_out_1_470;

    Conv_out_2[471]   <= conv_out_1_471;

    Conv_out_2[472]   <= conv_out_1_472;

    Conv_out_2[473]   <= conv_out_1_473;

    Conv_out_2[474]   <= conv_out_1_474;

    Conv_out_2[475]   <= conv_out_1_475;

    Conv_out_2[476]   <= conv_out_1_476;

    Conv_out_2[477]   <= conv_out_1_477;

    Conv_out_2[478]   <= conv_out_1_478;

    Conv_out_2[479]   <= conv_out_1_479;

    Conv_out_2[480]   <= conv_out_1_480;

    Conv_out_2[481]   <= conv_out_1_481;

    Conv_out_2[482]   <= conv_out_1_482;

    Conv_out_2[483]   <= conv_out_1_483;

    Conv_out_2[484]   <= conv_out_1_484;

    Conv_out_2[485]   <= conv_out_1_485;

    Conv_out_2[486]   <= conv_out_1_486;

    Conv_out_2[487]   <= conv_out_1_487;

    Conv_out_2[488]   <= conv_out_1_488;

    Conv_out_2[489]   <= conv_out_1_489;

    Conv_out_2[490]   <= conv_out_1_490;

    Conv_out_2[491]   <= conv_out_1_491;

    Conv_out_2[492]   <= conv_out_1_492;

    Conv_out_2[493]   <= conv_out_1_493;

    Conv_out_2[494]   <= conv_out_1_494;

    Conv_out_2[495]   <= conv_out_1_495;

    Conv_out_2[496]   <= conv_out_1_496;

    Conv_out_2[497]   <= conv_out_1_497;

    Conv_out_2[498]   <= conv_out_1_498;

    Conv_out_2[499]   <= conv_out_1_499;

    Conv_out_2[500]   <= conv_out_1_500;

    Conv_out_2[501]   <= conv_out_1_501;

    Conv_out_2[502]   <= conv_out_1_502;

    Conv_out_2[503]   <= conv_out_1_503;

    Conv_out_2[504]   <= conv_out_1_504;

    Conv_out_2[505]   <= conv_out_1_505;

    Conv_out_2[506]   <= conv_out_1_506;

    Conv_out_2[507]   <= conv_out_1_507;

    Conv_out_2[508]   <= conv_out_1_508;

    Conv_out_2[509]   <= conv_out_1_509;

    Conv_out_2[510]   <= conv_out_1_510;

    Conv_out_2[511]   <= conv_out_1_511;

    Conv_out_2[512]   <= conv_out_1_512;

    Conv_out_2[513]   <= conv_out_1_513;

    Conv_out_2[514]   <= conv_out_1_514;

    Conv_out_2[515]   <= conv_out_1_515;

    Conv_out_2[516]   <= conv_out_1_516;

    Conv_out_2[517]   <= conv_out_1_517;

    Conv_out_2[518]   <= conv_out_1_518;

    Conv_out_2[519]   <= conv_out_1_519;

    Conv_out_2[520]   <= conv_out_1_520;

    Conv_out_2[521]   <= conv_out_1_521;

    Conv_out_2[522]   <= conv_out_1_522;

    Conv_out_2[523]   <= conv_out_1_523;

    Conv_out_2[524]   <= conv_out_1_524;

    Conv_out_2[525]   <= conv_out_1_525;

    Conv_out_2[526]   <= conv_out_1_526;

    Conv_out_2[527]   <= conv_out_1_527;

    Conv_out_2[528]   <= conv_out_1_528;

    Conv_out_2[529]   <= conv_out_1_529;

    Conv_out_2[530]   <= conv_out_1_530;

    Conv_out_2[531]   <= conv_out_1_531;

    Conv_out_2[532]   <= conv_out_1_532;

    Conv_out_2[533]   <= conv_out_1_533;

    Conv_out_2[534]   <= conv_out_1_534;

    Conv_out_2[535]   <= conv_out_1_535;

    Conv_out_2[536]   <= conv_out_1_536;

    Conv_out_2[537]   <= conv_out_1_537;

    Conv_out_2[538]   <= conv_out_1_538;

    Conv_out_2[539]   <= conv_out_1_539;

    Conv_out_2[540]   <= conv_out_1_540;

    Conv_out_2[541]   <= conv_out_1_541;

    Conv_out_2[542]   <= conv_out_1_542;

    Conv_out_2[543]   <= conv_out_1_543;

    Conv_out_2[544]   <= conv_out_1_544;

    Conv_out_2[545]   <= conv_out_1_545;

    Conv_out_2[546]   <= conv_out_1_546;

    Conv_out_2[547]   <= conv_out_1_547;

    Conv_out_2[548]   <= conv_out_1_548;

    Conv_out_2[549]   <= conv_out_1_549;

    Conv_out_2[550]   <= conv_out_1_550;

    Conv_out_2[551]   <= conv_out_1_551;

    Conv_out_2[552]   <= conv_out_1_552;

    Conv_out_2[553]   <= conv_out_1_553;

    Conv_out_2[554]   <= conv_out_1_554;

    Conv_out_2[555]   <= conv_out_1_555;

    Conv_out_2[556]   <= conv_out_1_556;

    Conv_out_2[557]   <= conv_out_1_557;

    Conv_out_2[558]   <= conv_out_1_558;

    Conv_out_2[559]   <= conv_out_1_559;

    Conv_out_2[560]   <= conv_out_1_560;

    Conv_out_2[561]   <= conv_out_1_561;

    Conv_out_2[562]   <= conv_out_1_562;

    Conv_out_2[563]   <= conv_out_1_563;

    Conv_out_2[564]   <= conv_out_1_564;

    Conv_out_2[565]   <= conv_out_1_565;

    Conv_out_2[566]   <= conv_out_1_566;

    Conv_out_2[567]   <= conv_out_1_567;

    Conv_out_2[568]   <= conv_out_1_568;

    Conv_out_2[569]   <= conv_out_1_569;

    Conv_out_2[570]   <= conv_out_1_570;

    Conv_out_2[571]   <= conv_out_1_571;

    Conv_out_2[572]   <= conv_out_1_572;

    Conv_out_2[573]   <= conv_out_1_573;

    Conv_out_2[574]   <= conv_out_1_574;

    Conv_out_2[575]   <= conv_out_1_575;

    Conv_out_2[576]   <= conv_out_1_576;

    Conv_out_2[577]   <= conv_out_1_577;

    Conv_out_2[578]   <= conv_out_1_578;

    Conv_out_2[579]   <= conv_out_1_579;

    Conv_out_2[580]   <= conv_out_1_580;

    Conv_out_2[581]   <= conv_out_1_581;

    Conv_out_2[582]   <= conv_out_1_582;

    Conv_out_2[583]   <= conv_out_1_583;

    Conv_out_2[584]   <= conv_out_1_584;

    Conv_out_2[585]   <= conv_out_1_585;

    Conv_out_2[586]   <= conv_out_1_586;

    Conv_out_2[587]   <= conv_out_1_587;

    Conv_out_2[588]   <= conv_out_1_588;

    Conv_out_2[589]   <= conv_out_1_589;

    Conv_out_2[590]   <= conv_out_1_590;

    Conv_out_2[591]   <= conv_out_1_591;

    Conv_out_2[592]   <= conv_out_1_592;

    Conv_out_2[593]   <= conv_out_1_593;

    Conv_out_2[594]   <= conv_out_1_594;

    Conv_out_2[595]   <= conv_out_1_595;

    Conv_out_2[596]   <= conv_out_1_596;

    Conv_out_2[597]   <= conv_out_1_597;

    Conv_out_2[598]   <= conv_out_1_598;

    Conv_out_2[599]   <= conv_out_1_599;

    Conv_out_2[600]   <= conv_out_1_600;

    Conv_out_2[601]   <= conv_out_1_601;

    Conv_out_2[602]   <= conv_out_1_602;

    Conv_out_2[603]   <= conv_out_1_603;

    Conv_out_2[604]   <= conv_out_1_604;

    Conv_out_2[605]   <= conv_out_1_605;

    Conv_out_2[606]   <= conv_out_1_606;

    Conv_out_2[607]   <= conv_out_1_607;

    Conv_out_2[608]   <= conv_out_1_608;

    Conv_out_2[609]   <= conv_out_1_609;

    Conv_out_2[610]   <= conv_out_1_610;

    Conv_out_2[611]   <= conv_out_1_611;

    Conv_out_2[612]   <= conv_out_1_612;

    Conv_out_2[613]   <= conv_out_1_613;

    Conv_out_2[614]   <= conv_out_1_614;

    Conv_out_2[615]   <= conv_out_1_615;

    Conv_out_2[616]   <= conv_out_1_616;

    Conv_out_2[617]   <= conv_out_1_617;

    Conv_out_2[618]   <= conv_out_1_618;

    Conv_out_2[619]   <= conv_out_1_619;

    Conv_out_2[620]   <= conv_out_1_620;

    Conv_out_2[621]   <= conv_out_1_621;

    Conv_out_2[622]   <= conv_out_1_622;

    Conv_out_2[623]   <= conv_out_1_623;

    Conv_out_2[624]   <= conv_out_1_624;

    Conv_out_2[625]   <= conv_out_1_625;

    Conv_out_2[626]   <= conv_out_1_626;

    Conv_out_2[627]   <= conv_out_1_627;

    Conv_out_2[628]   <= conv_out_1_628;

    Conv_out_2[629]   <= conv_out_1_629;

    Conv_out_2[630]   <= conv_out_1_630;

    Conv_out_2[631]   <= conv_out_1_631;

    Conv_out_2[632]   <= conv_out_1_632;

    Conv_out_2[633]   <= conv_out_1_633;

    Conv_out_2[634]   <= conv_out_1_634;

    Conv_out_2[635]   <= conv_out_1_635;

    Conv_out_2[636]   <= conv_out_1_636;

    Conv_out_2[637]   <= conv_out_1_637;

    Conv_out_2[638]   <= conv_out_1_638;

    Conv_out_2[639]   <= conv_out_1_639;

    Conv_out_2[640]   <= conv_out_1_640;

    Conv_out_2[641]   <= conv_out_1_641;

    Conv_out_2[642]   <= conv_out_1_642;

    Conv_out_2[643]   <= conv_out_1_643;

    Conv_out_2[644]   <= conv_out_1_644;

    Conv_out_2[645]   <= conv_out_1_645;

    Conv_out_2[646]   <= conv_out_1_646;

    Conv_out_2[647]   <= conv_out_1_647;

    Conv_out_2[648]   <= conv_out_1_648;

    Conv_out_2[649]   <= conv_out_1_649;

    Conv_out_2[650]   <= conv_out_1_650;

    Conv_out_2[651]   <= conv_out_1_651;

    Conv_out_2[652]   <= conv_out_1_652;

    Conv_out_2[653]   <= conv_out_1_653;

    Conv_out_2[654]   <= conv_out_1_654;

    Conv_out_2[655]   <= conv_out_1_655;

    Conv_out_2[656]   <= conv_out_1_656;

    Conv_out_2[657]   <= conv_out_1_657;

    Conv_out_2[658]   <= conv_out_1_658;

    Conv_out_2[659]   <= conv_out_1_659;

    Conv_out_2[660]   <= conv_out_1_660;

    Conv_out_2[661]   <= conv_out_1_661;

    Conv_out_2[662]   <= conv_out_1_662;

    Conv_out_2[663]   <= conv_out_1_663;

    Conv_out_2[664]   <= conv_out_1_664;

    Conv_out_2[665]   <= conv_out_1_665;

    Conv_out_2[666]   <= conv_out_1_666;

    Conv_out_2[667]   <= conv_out_1_667;

    Conv_out_2[668]   <= conv_out_1_668;

    Conv_out_2[669]   <= conv_out_1_669;

    Conv_out_2[670]   <= conv_out_1_670;

    Conv_out_2[671]   <= conv_out_1_671;

    Conv_out_2[672]   <= conv_out_1_672;

    Conv_out_2[673]   <= conv_out_1_673;

    Conv_out_2[674]   <= conv_out_1_674;

    Conv_out_2[675]   <= conv_out_1_675;

    Conv_out_2[676]   <= conv_out_1_676;

    Conv_out_2[677]   <= conv_out_1_677;

    Conv_out_2[678]   <= conv_out_1_678;

    Conv_out_2[679]   <= conv_out_1_679;

    Conv_out_2[680]   <= conv_out_1_680;

    Conv_out_2[681]   <= conv_out_1_681;

    Conv_out_2[682]   <= conv_out_1_682;

    Conv_out_2[683]   <= conv_out_1_683;

    Conv_out_2[684]   <= conv_out_1_684;

    Conv_out_2[685]   <= conv_out_1_685;

    Conv_out_2[686]   <= conv_out_1_686;

    Conv_out_2[687]   <= conv_out_1_687;

    Conv_out_2[688]   <= conv_out_1_688;

    Conv_out_2[689]   <= conv_out_1_689;

    Conv_out_2[690]   <= conv_out_1_690;

    Conv_out_2[691]   <= conv_out_1_691;

    Conv_out_2[692]   <= conv_out_1_692;

    Conv_out_2[693]   <= conv_out_1_693;

    Conv_out_2[694]   <= conv_out_1_694;

    Conv_out_2[695]   <= conv_out_1_695;

    Conv_out_2[696]   <= conv_out_1_696;

    Conv_out_2[697]   <= conv_out_1_697;

    Conv_out_2[698]   <= conv_out_1_698;

    Conv_out_2[699]   <= conv_out_1_699;

    Conv_out_2[700]   <= conv_out_1_700;

    Conv_out_2[701]   <= conv_out_1_701;

    Conv_out_2[702]   <= conv_out_1_702;

    Conv_out_2[703]   <= conv_out_1_703;

    Conv_out_2[704]   <= conv_out_1_704;

    Conv_out_2[705]   <= conv_out_1_705;

    Conv_out_2[706]   <= conv_out_1_706;

    Conv_out_2[707]   <= conv_out_1_707;

    Conv_out_2[708]   <= conv_out_1_708;

    Conv_out_2[709]   <= conv_out_1_709;

    Conv_out_2[710]   <= conv_out_1_710;

    Conv_out_2[711]   <= conv_out_1_711;

    Conv_out_2[712]   <= conv_out_1_712;

    Conv_out_2[713]   <= conv_out_1_713;

    Conv_out_2[714]   <= conv_out_1_714;

    Conv_out_2[715]   <= conv_out_1_715;

    Conv_out_2[716]   <= conv_out_1_716;

    Conv_out_2[717]   <= conv_out_1_717;

    Conv_out_2[718]   <= conv_out_1_718;

    Conv_out_2[719]   <= conv_out_1_719;

    Conv_out_2[720]   <= conv_out_1_720;

    Conv_out_2[721]   <= conv_out_1_721;

    Conv_out_2[722]   <= conv_out_1_722;

    Conv_out_2[723]   <= conv_out_1_723;

    Conv_out_2[724]   <= conv_out_1_724;

    Conv_out_2[725]   <= conv_out_1_725;

    Conv_out_2[726]   <= conv_out_1_726;

    Conv_out_2[727]   <= conv_out_1_727;

    Conv_out_2[728]   <= conv_out_1_728;

    Conv_out_2[729]   <= conv_out_1_729;

    Conv_out_2[730]   <= conv_out_1_730;

    Conv_out_2[731]   <= conv_out_1_731;

    Conv_out_2[732]   <= conv_out_1_732;

    Conv_out_2[733]   <= conv_out_1_733;

    Conv_out_2[734]   <= conv_out_1_734;

    Conv_out_2[735]   <= conv_out_1_735;

    Conv_out_2[736]   <= conv_out_1_736;

    Conv_out_2[737]   <= conv_out_1_737;

    Conv_out_2[738]   <= conv_out_1_738;

    Conv_out_2[739]   <= conv_out_1_739;

    Conv_out_2[740]   <= conv_out_1_740;

    Conv_out_2[741]   <= conv_out_1_741;

    Conv_out_2[742]   <= conv_out_1_742;

    Conv_out_2[743]   <= conv_out_1_743;

    Conv_out_2[744]   <= conv_out_1_744;

    Conv_out_2[745]   <= conv_out_1_745;

    Conv_out_2[746]   <= conv_out_1_746;

    Conv_out_2[747]   <= conv_out_1_747;

    Conv_out_2[748]   <= conv_out_1_748;

    Conv_out_2[749]   <= conv_out_1_749;

    Conv_out_2[750]   <= conv_out_1_750;

    Conv_out_2[751]   <= conv_out_1_751;

    Conv_out_2[752]   <= conv_out_1_752;

    Conv_out_2[753]   <= conv_out_1_753;

    Conv_out_2[754]   <= conv_out_1_754;

    Conv_out_2[755]   <= conv_out_1_755;

    Conv_out_2[756]   <= conv_out_1_756;

    Conv_out_2[757]   <= conv_out_1_757;

    Conv_out_2[758]   <= conv_out_1_758;

    Conv_out_2[759]   <= conv_out_1_759;

    Conv_out_2[760]   <= conv_out_1_760;

    Conv_out_2[761]   <= conv_out_1_761;

    Conv_out_2[762]   <= conv_out_1_762;

    Conv_out_2[763]   <= conv_out_1_763;

    Conv_out_2[764]   <= conv_out_1_764;

    Conv_out_2[765]   <= conv_out_1_765;

    Conv_out_2[766]   <= conv_out_1_766;

    Conv_out_2[767]   <= conv_out_1_767;

    Conv_out_2[768]   <= conv_out_1_768;

    Conv_out_2[769]   <= conv_out_1_769;

    Conv_out_2[770]   <= conv_out_1_770;

    Conv_out_2[771]   <= conv_out_1_771;

    Conv_out_2[772]   <= conv_out_1_772;

    Conv_out_2[773]   <= conv_out_1_773;

    Conv_out_2[774]   <= conv_out_1_774;

    Conv_out_2[775]   <= conv_out_1_775;

    Conv_out_2[776]   <= conv_out_1_776;

    Conv_out_2[777]   <= conv_out_1_777;

    Conv_out_2[778]   <= conv_out_1_778;

    Conv_out_2[779]   <= conv_out_1_779;

    Conv_out_2[780]   <= conv_out_1_780;

    Conv_out_2[781]   <= conv_out_1_781;

    Conv_out_2[782]   <= conv_out_1_782;

    Conv_out_2[783]   <= conv_out_1_783;

end

//   integer file;

//   initial begin    
//        #5000;
//        file = $fopen("Conv_1.mem", "w"); 
//        $fdisplay(file, "%h", Conv_out);
//    end

    
endmodule
